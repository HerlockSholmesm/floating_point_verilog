module dp_sqrt(input [63:0]x, output reg[63:0] y);

reg[51:0]x_mantissa;
reg[10:0]x_exponent;
reg x_sign;
reg[51:0]y_mantissa;
reg[10:0]y_exponent;
reg y_sign;
//
reg[53:0]ix;
reg [26:0] r;
reg [26:0] q;
integer i;

always @(x)
begin
x_mantissa = x[51:0];
x_exponent = x[62:52];
x_sign = x[63];
y_sign = 1'b0;
//
r[26] = 1'b0;
q[26] = 1'b0;

if(x_exponent==11'b0000_0000_000)
begin
    y_exponent={1'b0,x_exponent[10:1]}+511;
//
    ix={1'b1,x_mantissa,2'b00};
    y_mantissa=52'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
else if (x_exponent==11'b11111111111)
begin
    y_exponent={1'b0,x_exponent[10:1]}+512;
    ix={2'b01,x_mantissa,1'b0};
    y_mantissa=52'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end
else
begin
    if(x_exponent[0]==1'b1)
    begin
        y_exponent={1'b0,x_exponent[10:1]}+512;
        ix={2'b01,x_mantissa,1'b0};
    end
    else
    begin
        y_exponent={1'b0,x_exponent[10:1]}+511;
        ix={1'b1,x_mantissa,2'b00};
    end
    
    y_mantissa=52'b0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
end

begin //loop
if (r[26:25+1] == 0)
 	 r[26:25] = ix[2*25+1:2*25] - 2'b01;
else 
 	 r[26:25] = ix[2*25+1:2*25] + 2'b11;
	 
if (r[26:25] == 0)
 	 q[26:25] = {q[26:25+1],1'b1};
 else
 	 q[26:25] = {q[26:25+1],1'b0};
#100;if (r[26] == 0)
 	 r[26:24] = { r[26:24+1], ix[2*24+1:2*24]} - {q[25:24+1],2'b01};
else 
 	 r[26:24] = { r[26:24+1], ix[2*24+1:2*24]} + {q[25:24+1],2'b11};
if (r[26] == 0)
 	 q[26:24] = {q[26:24+1],1'b1};
 else
 	 q[26:24] = {q[26:24+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:23] = { r[26:23+1], ix[2*23+1:2*23]} - {q[25:23+1],2'b01};
else 
 	 r[26:23] = { r[26:23+1], ix[2*23+1:2*23]} + {q[25:23+1],2'b11};
if (r[26] == 0)
 	 q[26:23] = {q[26:23+1],1'b1};
 else
 	 q[26:23] = {q[26:23+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:22] = { r[26:22+1], ix[2*22+1:2*22]} - {q[25:22+1],2'b01};
else 
 	 r[26:22] = { r[26:22+1], ix[2*22+1:2*22]} + {q[25:22+1],2'b11};
if (r[26] == 0)
 	 q[26:22] = {q[26:22+1],1'b1};
 else
 	 q[26:22] = {q[26:22+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:21] = { r[26:21+1], ix[2*21+1:2*21]} - {q[25:21+1],2'b01};
else 
 	 r[26:21] = { r[26:21+1], ix[2*21+1:2*21]} + {q[25:21+1],2'b11};
if (r[26] == 0)
 	 q[26:21] = {q[26:21+1],1'b1};
 else
 	 q[26:21] = {q[26:21+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:20] = { r[26:20+1], ix[2*20+1:2*20]} - {q[25:20+1],2'b01};
else 
 	 r[26:20] = { r[26:20+1], ix[2*20+1:2*20]} + {q[25:20+1],2'b11};
if (r[26] == 0)
 	 q[26:20] = {q[26:20+1],1'b1};
 else
 	 q[26:20] = {q[26:20+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:19] = { r[26:19+1], ix[2*19+1:2*19]} - {q[25:19+1],2'b01};
else 
 	 r[26:19] = { r[26:19+1], ix[2*19+1:2*19]} + {q[25:19+1],2'b11};
if (r[26] == 0)
 	 q[26:19] = {q[26:19+1],1'b1};
 else
 	 q[26:19] = {q[26:19+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:18] = { r[26:18+1], ix[2*18+1:2*18]} - {q[25:18+1],2'b01};
else 
 	 r[26:18] = { r[26:18+1], ix[2*18+1:2*18]} + {q[25:18+1],2'b11};
if (r[26] == 0)
 	 q[26:18] = {q[26:18+1],1'b1};
 else
 	 q[26:18] = {q[26:18+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:17] = { r[26:17+1], ix[2*17+1:2*17]} - {q[25:17+1],2'b01};
else 
 	 r[26:17] = { r[26:17+1], ix[2*17+1:2*17]} + {q[25:17+1],2'b11};
if (r[26] == 0)
 	 q[26:17] = {q[26:17+1],1'b1};
 else
 	 q[26:17] = {q[26:17+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:16] = { r[26:16+1], ix[2*16+1:2*16]} - {q[25:16+1],2'b01};
else 
 	 r[26:16] = { r[26:16+1], ix[2*16+1:2*16]} + {q[25:16+1],2'b11};
if (r[26] == 0)
 	 q[26:16] = {q[26:16+1],1'b1};
 else
 	 q[26:16] = {q[26:16+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:15] = { r[26:15+1], ix[2*15+1:2*15]} - {q[25:15+1],2'b01};
else 
 	 r[26:15] = { r[26:15+1], ix[2*15+1:2*15]} + {q[25:15+1],2'b11};
if (r[26] == 0)
 	 q[26:15] = {q[26:15+1],1'b1};
 else
 	 q[26:15] = {q[26:15+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:14] = { r[26:14+1], ix[2*14+1:2*14]} - {q[25:14+1],2'b01};
else 
 	 r[26:14] = { r[26:14+1], ix[2*14+1:2*14]} + {q[25:14+1],2'b11};
if (r[26] == 0)
 	 q[26:14] = {q[26:14+1],1'b1};
 else
 	 q[26:14] = {q[26:14+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:13] = { r[26:13+1], ix[2*13+1:2*13]} - {q[25:13+1],2'b01};
else 
 	 r[26:13] = { r[26:13+1], ix[2*13+1:2*13]} + {q[25:13+1],2'b11};
if (r[26] == 0)
 	 q[26:13] = {q[26:13+1],1'b1};
 else
 	 q[26:13] = {q[26:13+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:12] = { r[26:12+1], ix[2*12+1:2*12]} - {q[25:12+1],2'b01};
else 
 	 r[26:12] = { r[26:12+1], ix[2*12+1:2*12]} + {q[25:12+1],2'b11};
if (r[26] == 0)
 	 q[26:12] = {q[26:12+1],1'b1};
 else
 	 q[26:12] = {q[26:12+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:11] = { r[26:11+1], ix[2*11+1:2*11]} - {q[25:11+1],2'b01};
else 
 	 r[26:11] = { r[26:11+1], ix[2*11+1:2*11]} + {q[25:11+1],2'b11};
if (r[26] == 0)
 	 q[26:11] = {q[26:11+1],1'b1};
 else
 	 q[26:11] = {q[26:11+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:10] = { r[26:10+1], ix[2*10+1:2*10]} - {q[25:10+1],2'b01};
else 
 	 r[26:10] = { r[26:10+1], ix[2*10+1:2*10]} + {q[25:10+1],2'b11};
if (r[26] == 0)
 	 q[26:10] = {q[26:10+1],1'b1};
 else
 	 q[26:10] = {q[26:10+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:9] = { r[26:9+1], ix[2*9+1:2*9]} - {q[25:9+1],2'b01};
else 
 	 r[26:9] = { r[26:9+1], ix[2*9+1:2*9]} + {q[25:9+1],2'b11};
if (r[26] == 0)
 	 q[26:9] = {q[26:9+1],1'b1};
 else
 	 q[26:9] = {q[26:9+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:8] = { r[26:8+1], ix[2*8+1:2*8]} - {q[25:8+1],2'b01};
else 
 	 r[26:8] = { r[26:8+1], ix[2*8+1:2*8]} + {q[25:8+1],2'b11};
if (r[26] == 0)
 	 q[26:8] = {q[26:8+1],1'b1};
 else
 	 q[26:8] = {q[26:8+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:7] = { r[26:7+1], ix[2*7+1:2*7]} - {q[25:7+1],2'b01};
else 
 	 r[26:7] = { r[26:7+1], ix[2*7+1:2*7]} + {q[25:7+1],2'b11};
if (r[26] == 0)
 	 q[26:7] = {q[26:7+1],1'b1};
 else
 	 q[26:7] = {q[26:7+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:6] = { r[26:6+1], ix[2*6+1:2*6]} - {q[25:6+1],2'b01};
else 
 	 r[26:6] = { r[26:6+1], ix[2*6+1:2*6]} + {q[25:6+1],2'b11};
if (r[26] == 0)
 	 q[26:6] = {q[26:6+1],1'b1};
 else
 	 q[26:6] = {q[26:6+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:5] = { r[26:5+1], ix[2*5+1:2*5]} - {q[25:5+1],2'b01};
else 
 	 r[26:5] = { r[26:5+1], ix[2*5+1:2*5]} + {q[25:5+1],2'b11};
if (r[26] == 0)
 	 q[26:5] = {q[26:5+1],1'b1};
 else
 	 q[26:5] = {q[26:5+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:4] = { r[26:4+1], ix[2*4+1:2*4]} - {q[25:4+1],2'b01};
else 
 	 r[26:4] = { r[26:4+1], ix[2*4+1:2*4]} + {q[25:4+1],2'b11};
if (r[26] == 0)
 	 q[26:4] = {q[26:4+1],1'b1};
 else
 	 q[26:4] = {q[26:4+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:3] = { r[26:3+1], ix[2*3+1:2*3]} - {q[25:3+1],2'b01};
else 
 	 r[26:3] = { r[26:3+1], ix[2*3+1:2*3]} + {q[25:3+1],2'b11};
if (r[26] == 0)
 	 q[26:3] = {q[26:3+1],1'b1};
 else
 	 q[26:3] = {q[26:3+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:2] = { r[26:2+1], ix[2*2+1:2*2]} - {q[25:2+1],2'b01};
else 
 	 r[26:2] = { r[26:2+1], ix[2*2+1:2*2]} + {q[25:2+1],2'b11};
if (r[26] == 0)
 	 q[26:2] = {q[26:2+1],1'b1};
 else
 	 q[26:2] = {q[26:2+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:1] = { r[26:1+1], ix[2*1+1:2*1]} - {q[25:1+1],2'b01};
else 
 	 r[26:1] = { r[26:1+1], ix[2*1+1:2*1]} + {q[25:1+1],2'b11};
if (r[26] == 0)
 	 q[26:1] = {q[26:1+1],1'b1};
 else
 	 q[26:1] = {q[26:1+1],1'b0};
#100;

if (r[26] == 0)
 	 r[26:0] = { r[26:0+1], ix[2*0+1:2*0]} - {q[25:0+1],2'b01};
else 
 	 r[26:0] = { r[26:0+1], ix[2*0+1:2*0]} + {q[25:0+1],2'b11};
if (r[26] == 0)
 	 q[26:0] = {q[26:0+1],1'b1};
 else
 	 q[26:0] = {q[26:0+1],1'b0};
#100;







end

if (r[26] == 0) 
	r[26:0] = r[26:0] + {q[25:0],1'b1};


//
begin    
y_mantissa = {10'b0000_0000_00, q[12:0]};	
y[51:0]=y_mantissa;
y[62:52]=y_exponent;
y[63]=y_sign;
end
end
endmodule

