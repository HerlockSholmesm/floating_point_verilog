module sp_sqrt(input [31:0]x, output reg[31:0] y);

reg[22:0]x_mantissa;
reg[7:0]x_exponent;
reg x_sign;
reg[22:0]y_mantissa;
reg[7:0]y_exponent;
reg y_sign;
reg[25:0]ix;
reg [12:0] r;
reg [12:0] q;
integer i;

always @(x)
begin
x_mantissa = x[22:0];
x_exponent = x[30:23];
x_sign = x[31];
y_sign = 1'b0;
r[12] = 1'b0;
q[12] = 1'b0;

if(x_exponent==8'b00000000)
begin
    y_exponent={1'b0,x_exponent[7:1]}+63;
    ix={1'b0,x_mantissa,2'b00};
    y_mantissa=23'b0000_0000_0000_0000_0000_000;
end
else if (x_exponent==8'b11111111)
begin
    y_exponent={1'b0,x_exponent[7:1]}+64;
    ix={2'b00,x_mantissa,1'b0};
    y_mantissa=23'b0000_0000_0000_0000_0000_000;
end
else
begin
    if(x_exponent[0]==1'b1)
    begin
        y_exponent={1'b0,x_exponent[7:1]}+64;
        ix={2'b01,x_mantissa,1'b0};
    end
    else
    begin
        y_exponent={1'b0,x_exponent[7:1]}+63;
        ix={1'b1,x_mantissa,2'b00};
    end
    
    y_mantissa=23'b0000_0000_0000_0000_0000_000;
end
///after trying to model with clk I failed. so I tried to do it with loop.
begin //loop
if (r[12] == 0)
 	 r[12:11] = ix[2*11+1:2*11] - 2'b01;
else 
 	 r[12:11] = ix[2*11+1:2*11] + 2'b11;
	 
if (r[12] == 0)
 	 q[12:11] = {q[12:11+1],1'b1};
 else
 	 q[12:11] = {q[12:11+1],1'b0};
#100;
if (r[12] == 0)
 	 r[12:10] = { r[11:10+1], ix[2*10+1:2*10]} - {q[11:10+1],2'b01};
else 
 	 r[12:10] = { r[11:10+1], ix[2*10+1:2*10]} + {q[11:10+1],2'b11};
if (r[12] == 0)
 	 q[12:10] = {q[12:10+1],1'b1};
 else
 	 q[12:10] = {q[12:10+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:9] = { r[11:9+1], ix[2*9+1:2*9]} - {q[11:9+1],2'b01};
else 
 	 r[12:9] = { r[11:9+1], ix[2*9+1:2*9]} + {q[11:9+1],2'b11};
if (r[12] == 0)
 	 q[12:9] = {q[12:9+1],1'b1};
 else
 	 q[12:9] = {q[12:9+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:8] = { r[11:8+1], ix[2*8+1:2*8]} - {q[11:8+1],2'b01};
else 
 	 r[12:8] = { r[11:8+1], ix[2*8+1:2*8]} + {q[11:8+1],2'b11};
if (r[12] == 0)
 	 q[12:8] = {q[12:8+1],1'b1};
 else
 	 q[12:8] = {q[12:8+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:7] = { r[11:7+1], ix[2*7+1:2*7]} - {q[11:7+1],2'b01};
else 
 	 r[12:7] = { r[11:7+1], ix[2*7+1:2*7]} + {q[11:7+1],2'b11};
if (r[12] == 0)
 	 q[12:7] = {q[12:7+1],1'b1};
 else
 	 q[12:7] = {q[12:7+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:6] = { r[11:6+1], ix[2*6+1:2*6]} - {q[11:6+1],2'b01};
else 
 	 r[12:6] = { r[11:6+1], ix[2*6+1:2*6]} + {q[11:6+1],2'b11};
if (r[12] == 0)
 	 q[12:6] = {q[12:6+1],1'b1};
 else
 	 q[12:6] = {q[12:6+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:5] = { r[11:5+1], ix[2*5+1:2*5]} - {q[11:5+1],2'b01};
else 
 	 r[12:5] = { r[11:5+1], ix[2*5+1:2*5]} + {q[11:5+1],2'b11};
if (r[12] == 0)
 	 q[12:5] = {q[12:5+1],1'b1};
 else
 	 q[12:5] = {q[12:5+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:4] = { r[11:4+1], ix[2*4+1:2*4]} - {q[11:4+1],2'b01};
else 
 	 r[12:4] = { r[11:4+1], ix[2*4+1:2*4]} + {q[11:4+1],2'b11};
if (r[12] == 0)
 	 q[12:4] = {q[12:4+1],1'b1};
 else
 	 q[12:4] = {q[12:4+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:3] = { r[11:3+1], ix[2*3+1:2*3]} - {q[11:3+1],2'b01};
else 
 	 r[12:3] = { r[11:3+1], ix[2*3+1:2*3]} + {q[11:3+1],2'b11};
if (r[12] == 0)
 	 q[12:3] = {q[12:3+1],1'b1};
 else
 	 q[12:3] = {q[12:3+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:2] = { r[11:2+1], ix[2*2+1:2*2]} - {q[11:2+1],2'b01};
else 
 	 r[12:2] = { r[11:2+1], ix[2*2+1:2*2]} + {q[11:2+1],2'b11};
if (r[12] == 0)
 	 q[12:2] = {q[12:2+1],1'b1};
 else
 	 q[12:2] = {q[12:2+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:1] = { r[11:1+1], ix[2*1+1:2*1]} - {q[11:1+1],2'b01};
else 
 	 r[12:1] = { r[11:1+1], ix[2*1+1:2*1]} + {q[11:1+1],2'b11};
if (r[12] == 0)
 	 q[12:1] = {q[12:1+1],1'b1};
 else
 	 q[12:1] = {q[12:1+1],1'b0};
#100;

if (r[12] == 0)
 	 r[12:0] = { r[11:0+1], ix[2*0+1:2*0]} - {q[11:0+1],2'b01};
else 
 	 r[12:0] = { r[11:0+1], ix[2*0+1:2*0]} + {q[11:0+1],2'b11};
if (r[12] == 0)
 	 q[12:0] = {q[12:0+1],1'b1};
 else
 	 q[12:0] = {q[12:0+1],1'b0};
#100;




end

if (r[12:0] < 0) 
	r[12:0] = r[12:0] + {q[11:0],1'b1};

begin    
y_mantissa = {10'b0000_0000_00, q[12:0]};	
y[22:0]=y_mantissa;
y[30:23]=y_exponent;
y[31]=y_sign;
end
end
endmodule
