-- megafunction wizard: %ALTFP_SQRT%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_sqrt 

-- ============================================================
-- File Name: fp_sqrt_dp.vhd
-- Megafunction Name(s):
-- 			altfp_sqrt
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.0 Build 132 02/25/2009 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altfp_sqrt CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix II" PIPELINE=30 ROUNDING="TO_NEAREST" WIDTH_EXP=11 WIDTH_MAN=52 aclr clk_en clock data result
--VERSION_BEGIN 9.0 cbx_altfp_sqrt 2008:05:19:10:48:19:SJ cbx_cycloneii 2008:05:19:10:57:37:SJ cbx_lpm_add_sub 2008:12:09:22:11:50:SJ cbx_mgl 2009:01:29:16:12:07:SJ cbx_stratix 2008:09:18:16:08:35:SJ cbx_stratixii 2008:11:14:16:08:42:SJ  VERSION_END


--alt_sqrt_block CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Stratix II" PIPELINE=30 WIDTH_SQRT=54 aclr clken clock rad root_result
--VERSION_BEGIN 9.0 cbx_altfp_sqrt 2008:05:19:10:48:19:SJ cbx_cycloneii 2008:05:19:10:57:37:SJ cbx_lpm_add_sub 2008:12:09:22:11:50:SJ cbx_mgl 2009:01:29:16:12:07:SJ cbx_stratix 2008:09:18:16:08:35:SJ cbx_stratixii 2008:11:14:16:08:42:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 54 reg 2383 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fp_sqrt_dp_alt_sqrt_block_kgb IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 rad	:	IN  STD_LOGIC_VECTOR (54 DOWNTO 0);
		 root_result	:	OUT  STD_LOGIC_VECTOR (53 DOWNTO 0)
	 ); 
 END fp_sqrt_dp_alt_sqrt_block_kgb;

 ARCHITECTURE RTL OF fp_sqrt_dp_alt_sqrt_block_kgb IS

	 SIGNAL	 q_ff0c	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff10c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff12c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff14c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff16c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff18c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff20c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff22c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff24c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff26c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff28c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff2c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff30c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff32c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff34c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff36c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff38c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff40c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff42c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff44c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff46c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff48c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff4c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff50c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff52c	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff6c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 q_ff8c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rad_ff11c	:	STD_LOGIC_VECTOR(43 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff11c_w_lg_w_lg_w_q_range3587w3590w3591w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_lg_w_q_range3587w3588w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_lg_w_q_range3587w3590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_lg_w_lg_w_lg_w_q_range3587w3590w3591w3592w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_rad_ff11c_w_q_range3587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff13c	:	STD_LOGIC_VECTOR(41 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff13c_w_lg_w_lg_w_q_range3649w3652w3653w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_lg_w_q_range3649w3650w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_lg_w_q_range3649w3652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_lg_w_lg_w_lg_w_q_range3649w3652w3653w3654w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_rad_ff13c_w_q_range3649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff15c	:	STD_LOGIC_VECTOR(39 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff15c_w_lg_w_lg_w_q_range3711w3714w3715w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_lg_w_q_range3711w3712w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_lg_w_q_range3711w3714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_lg_w_lg_w_lg_w_q_range3711w3714w3715w3716w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_rad_ff15c_w_q_range3711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff17c	:	STD_LOGIC_VECTOR(37 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff17c_w_lg_w_lg_w_q_range3773w3776w3777w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_lg_w_q_range3773w3774w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_lg_w_q_range3773w3776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_lg_w_lg_w_lg_w_q_range3773w3776w3777w3778w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_rad_ff17c_w_q_range3773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff19c	:	STD_LOGIC_VECTOR(35 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff19c_w_lg_w_lg_w_q_range3835w3838w3839w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_lg_w_q_range3835w3836w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_lg_w_q_range3835w3838w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_lg_w_lg_w_lg_w_q_range3835w3838w3839w3840w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_rad_ff19c_w_q_range3835w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff1c	:	STD_LOGIC_VECTOR(53 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff1c_w_lg_w_lg_w_q_range3277w3280w3281w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_lg_w_q_range3277w3278w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_lg_w_q_range3277w3280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_lg_w_lg_w_lg_w_q_range3277w3280w3281w3282w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_rad_ff1c_w_q_range3277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff21c	:	STD_LOGIC_VECTOR(33 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff21c_w_lg_w_lg_w_q_range3897w3900w3901w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_lg_w_q_range3897w3898w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_lg_w_q_range3897w3900w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_lg_w_lg_w_lg_w_q_range3897w3900w3901w3902w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_rad_ff21c_w_q_range3897w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff23c	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff23c_w_lg_w_lg_w_q_range3959w3962w3963w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_lg_w_q_range3959w3960w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_lg_w_q_range3959w3962w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_lg_w_lg_w_lg_w_q_range3959w3962w3963w3964w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_rad_ff23c_w_q_range3959w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff25c	:	STD_LOGIC_VECTOR(29 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff25c_w_lg_w_lg_w_q_range4020w4023w4024w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_rad_ff25c_w_lg_w_q_range4020w4021w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_rad_ff25c_w_lg_w_q_range4020w4023w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff25c_w_lg_w_lg_w_lg_w_q_range4020w4023w4024w4025w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_rad_ff25c_w_q_range4020w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff27c	:	STD_LOGIC_VECTOR(27 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff27c_w_lg_w_lg_w_q_range4083w4086w4087w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_rad_ff27c_w_lg_w_q_range4083w4084w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_rad_ff27c_w_lg_w_q_range4083w4086w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff27c_w_lg_w_lg_w_lg_w_q_range4083w4086w4087w4088w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_rad_ff27c_w_q_range4083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff29c	:	STD_LOGIC_VECTOR(28 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff29c_w_lg_w_lg_w_q_range4160w4163w4164w	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_rad_ff29c_w_lg_w_q_range4160w4161w	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_rad_ff29c_w_lg_w_q_range4160w4163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff29c_w_lg_w_lg_w_lg_w_q_range4160w4163w4164w4165w	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_rad_ff29c_w_q_range4160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff31c	:	STD_LOGIC_VECTOR(30 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff31c_w_lg_w_lg_w_q_range4237w4240w4241w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_rad_ff31c_w_lg_w_q_range4237w4238w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_rad_ff31c_w_lg_w_q_range4237w4240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff31c_w_lg_w_lg_w_lg_w_q_range4237w4240w4241w4242w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_rad_ff31c_w_q_range4237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff33c	:	STD_LOGIC_VECTOR(32 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff33c_w_lg_w_lg_w_q_range4314w4317w4318w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_rad_ff33c_w_lg_w_q_range4314w4315w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_rad_ff33c_w_lg_w_q_range4314w4317w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff33c_w_lg_w_lg_w_lg_w_q_range4314w4317w4318w4319w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_rad_ff33c_w_q_range4314w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff35c	:	STD_LOGIC_VECTOR(34 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff35c_w_lg_w_lg_w_q_range4391w4394w4395w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_rad_ff35c_w_lg_w_q_range4391w4392w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_rad_ff35c_w_lg_w_q_range4391w4394w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff35c_w_lg_w_lg_w_lg_w_q_range4391w4394w4395w4396w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_rad_ff35c_w_q_range4391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff37c	:	STD_LOGIC_VECTOR(36 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff37c_w_lg_w_lg_w_q_range4468w4471w4472w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_rad_ff37c_w_lg_w_q_range4468w4469w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_rad_ff37c_w_lg_w_q_range4468w4471w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff37c_w_lg_w_lg_w_lg_w_q_range4468w4471w4472w4473w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_rad_ff37c_w_q_range4468w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff39c	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff39c_w_lg_w_lg_w_q_range4545w4548w4549w	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_rad_ff39c_w_lg_w_q_range4545w4546w	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_rad_ff39c_w_lg_w_q_range4545w4548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff39c_w_lg_w_lg_w_lg_w_q_range4545w4548w4549w4550w	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_rad_ff39c_w_q_range4545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff3c	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff3c_w_lg_w_lg_w_q_range3339w3342w3343w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_lg_w_q_range3339w3340w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_lg_w_q_range3339w3342w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_lg_w_lg_w_lg_w_q_range3339w3342w3343w3344w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_rad_ff3c_w_q_range3339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff41c	:	STD_LOGIC_VECTOR(40 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff41c_w_lg_w_lg_w_q_range4622w4625w4626w	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_rad_ff41c_w_lg_w_q_range4622w4623w	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_rad_ff41c_w_lg_w_q_range4622w4625w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff41c_w_lg_w_lg_w_lg_w_q_range4622w4625w4626w4627w	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_rad_ff41c_w_q_range4622w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff43c	:	STD_LOGIC_VECTOR(42 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff43c_w_lg_w_lg_w_q_range4699w4702w4703w	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_rad_ff43c_w_lg_w_q_range4699w4700w	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_rad_ff43c_w_lg_w_q_range4699w4702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff43c_w_lg_w_lg_w_lg_w_q_range4699w4702w4703w4704w	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_rad_ff43c_w_q_range4699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff45c	:	STD_LOGIC_VECTOR(44 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff45c_w_lg_w_lg_w_q_range4776w4779w4780w	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_rad_ff45c_w_lg_w_q_range4776w4777w	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_rad_ff45c_w_lg_w_q_range4776w4779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff45c_w_lg_w_lg_w_lg_w_q_range4776w4779w4780w4781w	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_rad_ff45c_w_q_range4776w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff47c	:	STD_LOGIC_VECTOR(46 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff47c_w_lg_w_lg_w_q_range4853w4856w4857w	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_rad_ff47c_w_lg_w_q_range4853w4854w	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_rad_ff47c_w_lg_w_q_range4853w4856w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff47c_w_lg_w_lg_w_lg_w_q_range4853w4856w4857w4858w	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_rad_ff47c_w_q_range4853w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff49c	:	STD_LOGIC_VECTOR(48 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff49c_w_lg_w_lg_w_q_range4930w4933w4934w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_rad_ff49c_w_lg_w_q_range4930w4931w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_rad_ff49c_w_lg_w_q_range4930w4933w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff49c_w_lg_w_lg_w_lg_w_q_range4930w4933w4934w4935w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_rad_ff49c_w_q_range4930w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff51c	:	STD_LOGIC_VECTOR(50 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff51c_w_lg_w_lg_w_q_range5007w5010w5011w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_rad_ff51c_w_lg_w_q_range5007w5008w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_rad_ff51c_w_lg_w_q_range5007w5010w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff51c_w_lg_w_lg_w_lg_w_q_range5007w5010w5011w5012w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_rad_ff51c_w_q_range5007w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff5c	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff5c_w_lg_w_lg_w_q_range3401w3404w3405w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_lg_w_q_range3401w3402w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_lg_w_q_range3401w3404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_lg_w_lg_w_lg_w_q_range3401w3404w3405w3406w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_rad_ff5c_w_q_range3401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff7c	:	STD_LOGIC_VECTOR(47 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff7c_w_lg_w_lg_w_q_range3463w3466w3467w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_lg_w_q_range3463w3464w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_lg_w_q_range3463w3466w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_lg_w_lg_w_lg_w_q_range3463w3466w3467w3468w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_rad_ff7c_w_q_range3463w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 rad_ff9c	:	STD_LOGIC_VECTOR(45 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_rad_ff9c_w_lg_w_lg_w_q_range3525w3528w3529w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_lg_w_q_range3525w3526w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_lg_w_q_range3525w3528w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_lg_w_lg_w_lg_w_q_range3525w3528w3529w3530w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_rad_ff9c_w_q_range3525w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_add_sub10_dataa	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub10_datab	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub10_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub11_dataa	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_add_sub11_datab	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_add_sub11_result	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_add_sub12_dataa	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub12_datab	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub12_result	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_add_sub13_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub13_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub13_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub14_dataa	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub14_datab	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub14_result	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_add_sub15_dataa	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub15_datab	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub15_result	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_add_sub16_dataa	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub16_datab	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub16_result	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_add_sub17_dataa	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub17_datab	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub17_result	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_add_sub18_dataa	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_add_sub18_datab	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_add_sub18_result	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_add_sub19_dataa	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub19_datab	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub19_result	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_add_sub20_dataa	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_add_sub20_datab	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_add_sub20_result	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_add_sub21_dataa	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_add_sub21_datab	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_add_sub21_result	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_add_sub22_dataa	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_add_sub22_datab	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_add_sub22_result	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_add_sub23_dataa	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_add_sub23_datab	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_add_sub23_result	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_add_sub24_dataa	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub24_datab	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub24_result	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_add_sub25_dataa	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_sub25_datab	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_sub25_result	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_add_sub26_dataa	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_add_sub26_datab	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_add_sub26_result	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_add_sub27_dataa	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_add_sub27_datab	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_add_sub27_result	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_add_sub28_dataa	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_sub28_datab	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_sub28_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_add_sub29_dataa	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub29_datab	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub29_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub30_dataa	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add_sub30_datab	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add_sub30_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add_sub31_dataa	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub31_datab	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub31_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub32_dataa	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub32_datab	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub32_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_add_sub33_dataa	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add_sub33_datab	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add_sub33_result	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_add_sub34_dataa	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_add_sub34_datab	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_add_sub34_result	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_add_sub35_dataa	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub35_datab	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub35_result	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_add_sub36_dataa	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub36_datab	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub36_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_add_sub37_dataa	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_add_sub37_datab	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_add_sub37_result	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_add_sub38_dataa	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_add_sub38_datab	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_add_sub38_result	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_add_sub39_dataa	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_add_sub39_datab	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_add_sub39_result	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_add_sub4_dataa	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_add_sub4_datab	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_add_sub4_result	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_add_sub40_dataa	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_add_sub40_datab	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_add_sub40_result	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_add_sub41_dataa	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_add_sub41_datab	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_add_sub41_result	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_add_sub42_dataa	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_add_sub42_datab	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_add_sub42_result	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_add_sub43_dataa	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add_sub43_datab	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add_sub43_result	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_add_sub44_dataa	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_add_sub44_datab	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_add_sub44_result	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_add_sub45_dataa	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_add_sub45_datab	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_add_sub45_result	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_add_sub46_dataa	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_add_sub46_datab	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_add_sub46_result	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_add_sub47_dataa	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_add_sub47_datab	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_add_sub47_result	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_add_sub48_dataa	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_add_sub48_datab	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_add_sub48_result	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_add_sub49_dataa	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_add_sub49_datab	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_add_sub49_result	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_add_sub5_dataa	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub5_datab	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub5_result	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_add_sub50_dataa	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_add_sub50_datab	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_add_sub50_result	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_add_sub51_dataa	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_add_sub51_datab	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_add_sub51_result	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_add_sub52_dataa	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_add_sub52_datab	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_add_sub52_result	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_add_sub53_dataa	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_add_sub53_datab	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_add_sub53_result	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_add_sub54_dataa	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_add_sub54_datab	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_add_sub54_result	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_add_sub55_dataa	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_add_sub55_datab	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_add_sub55_result	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_add_sub56_dataa	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_add_sub56_datab	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_add_sub56_result	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_add_sub57_dataa	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_add_sub57_datab	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_add_sub57_result	:	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  wire_add_sub6_dataa	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_datab	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub6_result	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_add_sub7_dataa	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub7_datab	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub7_result	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_add_sub8_dataa	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub8_datab	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub8_result	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_add_sub9_dataa	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub9_datab	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_add_sub9_result	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w10c_range783w784w3559w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w12c_range865w866w3621w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w14c_range947w948w3683w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w16c_range1029w1030w3745w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w18c_range1111w1112w3807w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w20c_range1193w1194w3869w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w22c_range1275w1276w3931w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w24c_range1357w1358w3993w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w26c_range1439w1440w4052w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w28c_range1520w1521w4125w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w2c_range455w456w3311w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w30c_range1600w1601w4202w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w32c_range1680w1681w4279w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w34c_range1760w1761w4356w	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w36c_range1840w1841w4433w	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w38c_range1920w1921w4510w	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w40c_range2000w2001w4587w	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w42c_range2080w2081w4664w	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w44c_range2160w2161w4741w	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w46c_range2240w2241w4818w	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w48c_range2320w2321w4895w	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w4c_range537w538w3373w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w50c_range2400w2401w4972w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w52c_range448w449w5050w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w6c_range619w620w3435w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w8c_range701w702w3497w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w3557w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w3619w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w3681w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w3743w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w3805w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w3867w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w3929w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w3991w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w4050w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w4123w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w3309w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w4200w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w4277w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w4354w	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w4431w	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w4508w	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w4585w	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w4662w	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w4739w	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w4816w	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w4893w	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w3371w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w4970w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w5048w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w3433w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w3495w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w784w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w11c_range787w788w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w866w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w13c_range869w870w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w948w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w15c_range951w952w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w1030w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w17c_range1033w1034w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w1112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w19c_range1115w1116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w1c_range367w368w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w1194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w21c_range1197w1198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w1276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w23c_range1279w1280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w1358w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w25c_range1361w1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w1440w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w27c_range1443w1444w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w1521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w29c_range1523w1524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w456w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w1601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w31c_range1603w1604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w1681w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w33c_range1683w1684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w1761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w35c_range1763w1764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w1841w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w37c_range1843w1844w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w1921w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w39c_range1923w1924w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w3c_range459w460w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w2001w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w41c_range2003w2004w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w2081w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w43c_range2083w2084w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w2161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w45c_range2163w2164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w2241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w47c_range2243w2244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w2321w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w49c_range2323w2324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w538w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w2401w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w51c_range2403w2404w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w449w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w53c_range452w453w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w5c_range541w542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w7c_range623w624w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_addnode_w9c_range705w706w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w10c_range3524w3527w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w11c_range3556w3558w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w12c_range3586w3589w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w13c_range3618w3620w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w14c_range3648w3651w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w15c_range3680w3682w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w16c_range3710w3713w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w17c_range3742w3744w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w18c_range3772w3775w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w19c_range3804w3806w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w20c_range3834w3837w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w21c_range3866w3868w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w22c_range3896w3899w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w23c_range3928w3930w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w24c_range3958w3961w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w25c_range3990w3992w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w26c_range4019w4022w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w27c_range4049w4051w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w28c_range4082w4085w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w29c_range4122w4124w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w2c_range3276w3279w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w30c_range4159w4162w	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w31c_range4199w4201w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w32c_range4236w4239w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w33c_range4276w4278w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w34c_range4313w4316w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w35c_range4353w4355w	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w36c_range4390w4393w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w37c_range4430w4432w	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w38c_range4467w4470w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w39c_range4507w4509w	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w3c_range3308w3310w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w40c_range4544w4547w	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w41c_range4584w4586w	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w42c_range4621w4624w	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w43c_range4661w4663w	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w44c_range4698w4701w	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w45c_range4738w4740w	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w46c_range4775w4778w	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w47c_range4815w4817w	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w48c_range4852w4855w	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w49c_range4892w4894w	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w4c_range3338w3341w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w50c_range4929w4932w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w51c_range4969w4971w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w52c_range5006w5009w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w53c_range5047w5049w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w5c_range3370w3372w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w6c_range3400w3403w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w7c_range3432w3434w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w8c_range3462w3465w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_lg_w_qlevel_w9c_range3494w3496w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3560w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3622w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3684w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3746w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3808w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3870w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3932w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3994w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4053w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4126w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3312w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4203w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4280w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4357w	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4434w	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4511w	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4588w	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4665w	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4742w	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4819w	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4896w	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3374w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w4973w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w5051w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3436w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w3498w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  addnode_w0c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w10c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w11c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w12c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w13c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w14c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w15c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w16c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w17c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w18c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w19c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w1c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w20c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w21c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w22c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w23c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w24c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w25c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w26c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w27c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w28c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w29c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w2c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w30c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w31c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w32c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w33c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w34c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w35c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w36c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w37c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w38c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w39c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w3c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w40c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w41c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w42c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w43c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w44c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w45c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w46c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w47c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w48c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w49c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w4c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w50c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w51c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w52c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w53c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w5c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w6c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w7c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w8c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  addnode_w9c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  qlevel_w0c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  qlevel_w10c :	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  qlevel_w11c :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  qlevel_w12c :	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  qlevel_w13c :	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  qlevel_w14c :	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  qlevel_w15c :	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  qlevel_w16c :	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  qlevel_w17c :	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  qlevel_w18c :	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  qlevel_w19c :	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  qlevel_w1c :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  qlevel_w20c :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  qlevel_w21c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  qlevel_w22c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  qlevel_w23c :	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  qlevel_w24c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  qlevel_w25c :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  qlevel_w26c :	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  qlevel_w27c :	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  qlevel_w28c :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  qlevel_w29c :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  qlevel_w2c :	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  qlevel_w30c :	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  qlevel_w31c :	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  qlevel_w32c :	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  qlevel_w33c :	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  qlevel_w34c :	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  qlevel_w35c :	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  qlevel_w36c :	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  qlevel_w37c :	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  qlevel_w38c :	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  qlevel_w39c :	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  qlevel_w3c :	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  qlevel_w40c :	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  qlevel_w41c :	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  qlevel_w42c :	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  qlevel_w43c :	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  qlevel_w44c :	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  qlevel_w45c :	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  qlevel_w46c :	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  qlevel_w47c :	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  qlevel_w48c :	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  qlevel_w49c :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  qlevel_w4c :	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  qlevel_w50c :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  qlevel_w51c :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  qlevel_w52c :	STD_LOGIC_VECTOR (54 DOWNTO 0);
	 SIGNAL  qlevel_w53c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  qlevel_w5c :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  qlevel_w6c :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  qlevel_w7c :	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 SIGNAL  qlevel_w8c :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  qlevel_w9c :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  slevel_w0c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w10c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w11c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w12c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w13c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w14c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w15c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w16c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w17c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w18c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w19c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w1c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w20c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w21c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w22c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w23c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w24c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w25c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w26c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w27c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w28c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w29c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w2c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w30c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w31c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w32c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w33c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w34c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w35c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w36c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w37c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w38c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w39c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w3c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w40c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w41c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w42c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w43c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w44c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w45c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w46c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w47c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w48c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w49c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w4c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w50c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w51c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w52c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w53c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w5c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w6c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w7c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w8c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  slevel_w9c :	STD_LOGIC_VECTOR (55 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w10c_range783w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w11c_range346w	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w11c_range787w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w12c_range865w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w13c_range347w	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w13c_range869w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w14c_range947w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w15c_range348w	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w15c_range951w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w16c_range1029w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w17c_range349w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w17c_range1033w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w18c_range1111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w19c_range350w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w19c_range1115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w1c_range341w	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w1c_range367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w20c_range1193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w21c_range351w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w21c_range1197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w22c_range1275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w23c_range352w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w23c_range1279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w24c_range1357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w25c_range353w	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w25c_range1361w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w26c_range1439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w27c_range354w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w27c_range1443w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w28c_range1520w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w29c_range355w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w29c_range1523w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w2c_range455w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w30c_range1600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w31c_range356w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w31c_range1603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w32c_range1680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w33c_range357w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w33c_range1683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w34c_range1760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w35c_range358w	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w35c_range1763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w36c_range1840w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w37c_range359w	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w37c_range1843w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w38c_range1920w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w39c_range360w	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w39c_range1923w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w3c_range342w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w3c_range459w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w40c_range2000w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w41c_range361w	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w41c_range2003w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w42c_range2080w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w43c_range362w	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w43c_range2083w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w44c_range2160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w45c_range363w	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w45c_range2163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w46c_range2240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w47c_range2243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w47c_range364w	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w48c_range2320w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w49c_range2323w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w49c_range365w	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w4c_range537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w50c_range2400w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w51c_range366w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w51c_range2403w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w52c_range448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w53c_range452w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w5c_range541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w5c_range343w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w6c_range619w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w7c_range623w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w7c_range344w	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w8c_range701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w9c_range345w	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_addnode_w9c_range705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w10c_range3524w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w11c_range3556w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w12c_range3586w	:	STD_LOGIC_VECTOR (12 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w13c_range3618w	:	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w14c_range3648w	:	STD_LOGIC_VECTOR (14 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w15c_range3680w	:	STD_LOGIC_VECTOR (15 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w16c_range3710w	:	STD_LOGIC_VECTOR (16 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w17c_range3742w	:	STD_LOGIC_VECTOR (17 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w18c_range3772w	:	STD_LOGIC_VECTOR (18 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w19c_range3804w	:	STD_LOGIC_VECTOR (19 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w20c_range3834w	:	STD_LOGIC_VECTOR (20 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w21c_range3866w	:	STD_LOGIC_VECTOR (21 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w22c_range3896w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w23c_range3928w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w24c_range3958w	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w25c_range3990w	:	STD_LOGIC_VECTOR (25 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w26c_range4019w	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w27c_range4049w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w28c_range4082w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w29c_range4122w	:	STD_LOGIC_VECTOR (28 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w2c_range3276w	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w30c_range4159w	:	STD_LOGIC_VECTOR (29 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w31c_range4199w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w32c_range4236w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w33c_range4276w	:	STD_LOGIC_VECTOR (32 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w34c_range4313w	:	STD_LOGIC_VECTOR (33 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w35c_range4353w	:	STD_LOGIC_VECTOR (34 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w36c_range4390w	:	STD_LOGIC_VECTOR (35 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w37c_range4430w	:	STD_LOGIC_VECTOR (36 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w38c_range4467w	:	STD_LOGIC_VECTOR (37 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w39c_range4507w	:	STD_LOGIC_VECTOR (38 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w3c_range3308w	:	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w40c_range4544w	:	STD_LOGIC_VECTOR (39 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w41c_range4584w	:	STD_LOGIC_VECTOR (40 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w42c_range4621w	:	STD_LOGIC_VECTOR (41 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w43c_range4661w	:	STD_LOGIC_VECTOR (42 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w44c_range4698w	:	STD_LOGIC_VECTOR (43 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w45c_range4738w	:	STD_LOGIC_VECTOR (44 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w46c_range4775w	:	STD_LOGIC_VECTOR (45 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w47c_range4815w	:	STD_LOGIC_VECTOR (46 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w48c_range4852w	:	STD_LOGIC_VECTOR (47 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w49c_range4892w	:	STD_LOGIC_VECTOR (48 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w4c_range3338w	:	STD_LOGIC_VECTOR (4 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w50c_range4929w	:	STD_LOGIC_VECTOR (49 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w51c_range4969w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w52c_range5006w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w53c_range5047w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w5c_range3370w	:	STD_LOGIC_VECTOR (5 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w6c_range3400w	:	STD_LOGIC_VECTOR (6 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w7c_range3432w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w8c_range3462w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_alt_sqrt_block2_w_qlevel_w9c_range3494w	:	STD_LOGIC_VECTOR (9 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	loop0 : FOR i IN 0 TO 11 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w10c_range783w784w3559w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w784w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w11c_range3556w3558w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 13 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w12c_range865w866w3621w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w866w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w13c_range3618w3620w(i);
	END GENERATE loop1;
	loop2 : FOR i IN 0 TO 15 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w14c_range947w948w3683w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w948w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w15c_range3680w3682w(i);
	END GENERATE loop2;
	loop3 : FOR i IN 0 TO 17 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w16c_range1029w1030w3745w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w1030w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w17c_range3742w3744w(i);
	END GENERATE loop3;
	loop4 : FOR i IN 0 TO 19 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w18c_range1111w1112w3807w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w1112w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w19c_range3804w3806w(i);
	END GENERATE loop4;
	loop5 : FOR i IN 0 TO 21 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w20c_range1193w1194w3869w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w1194w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w21c_range3866w3868w(i);
	END GENERATE loop5;
	loop6 : FOR i IN 0 TO 23 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w22c_range1275w1276w3931w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w1276w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w23c_range3928w3930w(i);
	END GENERATE loop6;
	loop7 : FOR i IN 0 TO 25 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w24c_range1357w1358w3993w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w1358w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w25c_range3990w3992w(i);
	END GENERATE loop7;
	loop8 : FOR i IN 0 TO 27 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w26c_range1439w1440w4052w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w1440w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w27c_range4049w4051w(i);
	END GENERATE loop8;
	loop9 : FOR i IN 0 TO 28 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w28c_range1520w1521w4125w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w1521w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w29c_range4122w4124w(i);
	END GENERATE loop9;
	loop10 : FOR i IN 0 TO 3 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w2c_range455w456w3311w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w456w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w3c_range3308w3310w(i);
	END GENERATE loop10;
	loop11 : FOR i IN 0 TO 30 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w30c_range1600w1601w4202w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w1601w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w31c_range4199w4201w(i);
	END GENERATE loop11;
	loop12 : FOR i IN 0 TO 32 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w32c_range1680w1681w4279w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w1681w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w33c_range4276w4278w(i);
	END GENERATE loop12;
	loop13 : FOR i IN 0 TO 34 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w34c_range1760w1761w4356w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w1761w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w35c_range4353w4355w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 36 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w36c_range1840w1841w4433w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w1841w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w37c_range4430w4432w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 38 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w38c_range1920w1921w4510w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w1921w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w39c_range4507w4509w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 40 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w40c_range2000w2001w4587w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w2001w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w41c_range4584w4586w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 42 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w42c_range2080w2081w4664w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w2081w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w43c_range4661w4663w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 44 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w44c_range2160w2161w4741w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w2161w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w45c_range4738w4740w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 46 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w46c_range2240w2241w4818w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w2241w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w47c_range4815w4817w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 48 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w48c_range2320w2321w4895w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w2321w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w49c_range4892w4894w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 5 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w4c_range537w538w3373w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w538w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w5c_range3370w3372w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w50c_range2400w2401w4972w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w2401w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w51c_range4969w4971w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w52c_range448w449w5050w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w449w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w53c_range5047w5049w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 7 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w6c_range619w620w3435w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w620w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w7c_range3432w3434w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 9 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w8c_range701w702w3497w(i) <= wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w702w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w9c_range3494w3496w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 11 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w3557w(i) <= wire_alt_sqrt_block2_w_addnode_w10c_range783w(0) AND wire_alt_sqrt_block2_w_qlevel_w11c_range3556w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 13 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w3619w(i) <= wire_alt_sqrt_block2_w_addnode_w12c_range865w(0) AND wire_alt_sqrt_block2_w_qlevel_w13c_range3618w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 15 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w3681w(i) <= wire_alt_sqrt_block2_w_addnode_w14c_range947w(0) AND wire_alt_sqrt_block2_w_qlevel_w15c_range3680w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 17 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w3743w(i) <= wire_alt_sqrt_block2_w_addnode_w16c_range1029w(0) AND wire_alt_sqrt_block2_w_qlevel_w17c_range3742w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 19 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w3805w(i) <= wire_alt_sqrt_block2_w_addnode_w18c_range1111w(0) AND wire_alt_sqrt_block2_w_qlevel_w19c_range3804w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 21 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w3867w(i) <= wire_alt_sqrt_block2_w_addnode_w20c_range1193w(0) AND wire_alt_sqrt_block2_w_qlevel_w21c_range3866w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 23 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w3929w(i) <= wire_alt_sqrt_block2_w_addnode_w22c_range1275w(0) AND wire_alt_sqrt_block2_w_qlevel_w23c_range3928w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 25 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w3991w(i) <= wire_alt_sqrt_block2_w_addnode_w24c_range1357w(0) AND wire_alt_sqrt_block2_w_qlevel_w25c_range3990w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 27 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w4050w(i) <= wire_alt_sqrt_block2_w_addnode_w26c_range1439w(0) AND wire_alt_sqrt_block2_w_qlevel_w27c_range4049w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 28 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w4123w(i) <= wire_alt_sqrt_block2_w_addnode_w28c_range1520w(0) AND wire_alt_sqrt_block2_w_qlevel_w29c_range4122w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 3 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w3309w(i) <= wire_alt_sqrt_block2_w_addnode_w2c_range455w(0) AND wire_alt_sqrt_block2_w_qlevel_w3c_range3308w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 30 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w4200w(i) <= wire_alt_sqrt_block2_w_addnode_w30c_range1600w(0) AND wire_alt_sqrt_block2_w_qlevel_w31c_range4199w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 32 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w4277w(i) <= wire_alt_sqrt_block2_w_addnode_w32c_range1680w(0) AND wire_alt_sqrt_block2_w_qlevel_w33c_range4276w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 34 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w4354w(i) <= wire_alt_sqrt_block2_w_addnode_w34c_range1760w(0) AND wire_alt_sqrt_block2_w_qlevel_w35c_range4353w(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 36 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w4431w(i) <= wire_alt_sqrt_block2_w_addnode_w36c_range1840w(0) AND wire_alt_sqrt_block2_w_qlevel_w37c_range4430w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 38 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w4508w(i) <= wire_alt_sqrt_block2_w_addnode_w38c_range1920w(0) AND wire_alt_sqrt_block2_w_qlevel_w39c_range4507w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 40 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w4585w(i) <= wire_alt_sqrt_block2_w_addnode_w40c_range2000w(0) AND wire_alt_sqrt_block2_w_qlevel_w41c_range4584w(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 42 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w4662w(i) <= wire_alt_sqrt_block2_w_addnode_w42c_range2080w(0) AND wire_alt_sqrt_block2_w_qlevel_w43c_range4661w(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 44 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w4739w(i) <= wire_alt_sqrt_block2_w_addnode_w44c_range2160w(0) AND wire_alt_sqrt_block2_w_qlevel_w45c_range4738w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 46 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w4816w(i) <= wire_alt_sqrt_block2_w_addnode_w46c_range2240w(0) AND wire_alt_sqrt_block2_w_qlevel_w47c_range4815w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 48 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w4893w(i) <= wire_alt_sqrt_block2_w_addnode_w48c_range2320w(0) AND wire_alt_sqrt_block2_w_qlevel_w49c_range4892w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 5 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w3371w(i) <= wire_alt_sqrt_block2_w_addnode_w4c_range537w(0) AND wire_alt_sqrt_block2_w_qlevel_w5c_range3370w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w4970w(i) <= wire_alt_sqrt_block2_w_addnode_w50c_range2400w(0) AND wire_alt_sqrt_block2_w_qlevel_w51c_range4969w(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w5048w(i) <= wire_alt_sqrt_block2_w_addnode_w52c_range448w(0) AND wire_alt_sqrt_block2_w_qlevel_w53c_range5047w(i);
	END GENERATE loop49;
	loop50 : FOR i IN 0 TO 7 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w3433w(i) <= wire_alt_sqrt_block2_w_addnode_w6c_range619w(0) AND wire_alt_sqrt_block2_w_qlevel_w7c_range3432w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 9 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w3495w(i) <= wire_alt_sqrt_block2_w_addnode_w8c_range701w(0) AND wire_alt_sqrt_block2_w_qlevel_w9c_range3494w(i);
	END GENERATE loop51;
	wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w784w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w10c_range783w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w11c_range787w788w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w11c_range787w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w866w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w12c_range865w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w13c_range869w870w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w13c_range869w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w948w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w14c_range947w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w15c_range951w952w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w15c_range951w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w1030w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w16c_range1029w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w17c_range1033w1034w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w17c_range1033w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w1112w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w18c_range1111w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w19c_range1115w1116w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w19c_range1115w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w1c_range367w368w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w1c_range367w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w1194w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w20c_range1193w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w21c_range1197w1198w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w21c_range1197w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w1276w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w22c_range1275w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w23c_range1279w1280w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w23c_range1279w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w1358w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w24c_range1357w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w25c_range1361w1362w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w25c_range1361w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w1440w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w26c_range1439w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w27c_range1443w1444w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w27c_range1443w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w1521w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w28c_range1520w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w29c_range1523w1524w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w29c_range1523w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w456w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w2c_range455w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w1601w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w30c_range1600w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w31c_range1603w1604w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w31c_range1603w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w1681w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w32c_range1680w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w33c_range1683w1684w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w33c_range1683w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w1761w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w34c_range1760w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w35c_range1763w1764w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w35c_range1763w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w1841w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w36c_range1840w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w37c_range1843w1844w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w37c_range1843w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w1921w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w38c_range1920w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w39c_range1923w1924w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w39c_range1923w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w3c_range459w460w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w3c_range459w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w2001w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w40c_range2000w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w41c_range2003w2004w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w41c_range2003w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w2081w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w42c_range2080w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w43c_range2083w2084w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w43c_range2083w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w2161w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w44c_range2160w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w45c_range2163w2164w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w45c_range2163w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w2241w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w46c_range2240w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w47c_range2243w2244w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w47c_range2243w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w2321w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w48c_range2320w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w49c_range2323w2324w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w49c_range2323w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w538w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w4c_range537w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w2401w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w50c_range2400w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w51c_range2403w2404w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w51c_range2403w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w449w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w52c_range448w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w53c_range452w453w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w53c_range452w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w5c_range541w542w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w5c_range541w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w620w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w6c_range619w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w7c_range623w624w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w7c_range623w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w702w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w8c_range701w(0);
	wire_alt_sqrt_block2_w_lg_w_addnode_w9c_range705w706w(0) <= NOT wire_alt_sqrt_block2_w_addnode_w9c_range705w(0);
	loop52 : FOR i IN 0 TO 10 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w10c_range3524w3527w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w10c_range3524w(i);
	END GENERATE loop52;
	loop53 : FOR i IN 0 TO 11 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w11c_range3556w3558w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w11c_range3556w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 12 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w12c_range3586w3589w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w12c_range3586w(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 13 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w13c_range3618w3620w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w13c_range3618w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 14 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w14c_range3648w3651w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w14c_range3648w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 15 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w15c_range3680w3682w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w15c_range3680w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 16 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w16c_range3710w3713w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w16c_range3710w(i);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 17 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w17c_range3742w3744w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w17c_range3742w(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 18 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w18c_range3772w3775w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w18c_range3772w(i);
	END GENERATE loop60;
	loop61 : FOR i IN 0 TO 19 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w19c_range3804w3806w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w19c_range3804w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 20 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w20c_range3834w3837w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w20c_range3834w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 21 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w21c_range3866w3868w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w21c_range3866w(i);
	END GENERATE loop63;
	loop64 : FOR i IN 0 TO 22 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w22c_range3896w3899w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w22c_range3896w(i);
	END GENERATE loop64;
	loop65 : FOR i IN 0 TO 23 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w23c_range3928w3930w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w23c_range3928w(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 24 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w24c_range3958w3961w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w24c_range3958w(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 25 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w25c_range3990w3992w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w25c_range3990w(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 26 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w26c_range4019w4022w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w26c_range4019w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 27 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w27c_range4049w4051w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w27c_range4049w(i);
	END GENERATE loop69;
	loop70 : FOR i IN 0 TO 27 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w28c_range4082w4085w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w28c_range4082w(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 28 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w29c_range4122w4124w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w29c_range4122w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 2 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w2c_range3276w3279w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w2c_range3276w(i);
	END GENERATE loop72;
	loop73 : FOR i IN 0 TO 29 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w30c_range4159w4162w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w30c_range4159w(i);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 30 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w31c_range4199w4201w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w31c_range4199w(i);
	END GENERATE loop74;
	loop75 : FOR i IN 0 TO 31 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w32c_range4236w4239w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w32c_range4236w(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 32 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w33c_range4276w4278w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w33c_range4276w(i);
	END GENERATE loop76;
	loop77 : FOR i IN 0 TO 33 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w34c_range4313w4316w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w34c_range4313w(i);
	END GENERATE loop77;
	loop78 : FOR i IN 0 TO 34 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w35c_range4353w4355w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w35c_range4353w(i);
	END GENERATE loop78;
	loop79 : FOR i IN 0 TO 35 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w36c_range4390w4393w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w36c_range4390w(i);
	END GENERATE loop79;
	loop80 : FOR i IN 0 TO 36 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w37c_range4430w4432w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w37c_range4430w(i);
	END GENERATE loop80;
	loop81 : FOR i IN 0 TO 37 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w38c_range4467w4470w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w38c_range4467w(i);
	END GENERATE loop81;
	loop82 : FOR i IN 0 TO 38 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w39c_range4507w4509w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w39c_range4507w(i);
	END GENERATE loop82;
	loop83 : FOR i IN 0 TO 3 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w3c_range3308w3310w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w3c_range3308w(i);
	END GENERATE loop83;
	loop84 : FOR i IN 0 TO 39 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w40c_range4544w4547w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w40c_range4544w(i);
	END GENERATE loop84;
	loop85 : FOR i IN 0 TO 40 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w41c_range4584w4586w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w41c_range4584w(i);
	END GENERATE loop85;
	loop86 : FOR i IN 0 TO 41 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w42c_range4621w4624w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w42c_range4621w(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 42 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w43c_range4661w4663w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w43c_range4661w(i);
	END GENERATE loop87;
	loop88 : FOR i IN 0 TO 43 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w44c_range4698w4701w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w44c_range4698w(i);
	END GENERATE loop88;
	loop89 : FOR i IN 0 TO 44 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w45c_range4738w4740w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w45c_range4738w(i);
	END GENERATE loop89;
	loop90 : FOR i IN 0 TO 45 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w46c_range4775w4778w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w46c_range4775w(i);
	END GENERATE loop90;
	loop91 : FOR i IN 0 TO 46 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w47c_range4815w4817w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w47c_range4815w(i);
	END GENERATE loop91;
	loop92 : FOR i IN 0 TO 47 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w48c_range4852w4855w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w48c_range4852w(i);
	END GENERATE loop92;
	loop93 : FOR i IN 0 TO 48 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w49c_range4892w4894w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w49c_range4892w(i);
	END GENERATE loop93;
	loop94 : FOR i IN 0 TO 4 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w4c_range3338w3341w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w4c_range3338w(i);
	END GENERATE loop94;
	loop95 : FOR i IN 0 TO 49 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w50c_range4929w4932w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w50c_range4929w(i);
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w51c_range4969w4971w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w51c_range4969w(i);
	END GENERATE loop96;
	loop97 : FOR i IN 0 TO 51 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w52c_range5006w5009w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w52c_range5006w(i);
	END GENERATE loop97;
	loop98 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w53c_range5047w5049w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w53c_range5047w(i);
	END GENERATE loop98;
	loop99 : FOR i IN 0 TO 5 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w5c_range3370w3372w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w5c_range3370w(i);
	END GENERATE loop99;
	loop100 : FOR i IN 0 TO 6 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w6c_range3400w3403w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w6c_range3400w(i);
	END GENERATE loop100;
	loop101 : FOR i IN 0 TO 7 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w7c_range3432w3434w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w7c_range3432w(i);
	END GENERATE loop101;
	loop102 : FOR i IN 0 TO 8 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w8c_range3462w3465w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w8c_range3462w(i);
	END GENERATE loop102;
	loop103 : FOR i IN 0 TO 9 GENERATE 
		wire_alt_sqrt_block2_w_lg_w_qlevel_w9c_range3494w3496w(i) <= NOT wire_alt_sqrt_block2_w_qlevel_w9c_range3494w(i);
	END GENERATE loop103;
	loop104 : FOR i IN 0 TO 11 GENERATE 
		wire_alt_sqrt_block2_w3560w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w10c_range783w784w3559w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w3557w(i);
	END GENERATE loop104;
	loop105 : FOR i IN 0 TO 13 GENERATE 
		wire_alt_sqrt_block2_w3622w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w12c_range865w866w3621w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w3619w(i);
	END GENERATE loop105;
	loop106 : FOR i IN 0 TO 15 GENERATE 
		wire_alt_sqrt_block2_w3684w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w14c_range947w948w3683w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w3681w(i);
	END GENERATE loop106;
	loop107 : FOR i IN 0 TO 17 GENERATE 
		wire_alt_sqrt_block2_w3746w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w16c_range1029w1030w3745w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w3743w(i);
	END GENERATE loop107;
	loop108 : FOR i IN 0 TO 19 GENERATE 
		wire_alt_sqrt_block2_w3808w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w18c_range1111w1112w3807w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w3805w(i);
	END GENERATE loop108;
	loop109 : FOR i IN 0 TO 21 GENERATE 
		wire_alt_sqrt_block2_w3870w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w20c_range1193w1194w3869w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w3867w(i);
	END GENERATE loop109;
	loop110 : FOR i IN 0 TO 23 GENERATE 
		wire_alt_sqrt_block2_w3932w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w22c_range1275w1276w3931w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w3929w(i);
	END GENERATE loop110;
	loop111 : FOR i IN 0 TO 25 GENERATE 
		wire_alt_sqrt_block2_w3994w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w24c_range1357w1358w3993w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w3991w(i);
	END GENERATE loop111;
	loop112 : FOR i IN 0 TO 27 GENERATE 
		wire_alt_sqrt_block2_w4053w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w26c_range1439w1440w4052w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w4050w(i);
	END GENERATE loop112;
	loop113 : FOR i IN 0 TO 28 GENERATE 
		wire_alt_sqrt_block2_w4126w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w28c_range1520w1521w4125w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w4123w(i);
	END GENERATE loop113;
	loop114 : FOR i IN 0 TO 3 GENERATE 
		wire_alt_sqrt_block2_w3312w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w2c_range455w456w3311w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w3309w(i);
	END GENERATE loop114;
	loop115 : FOR i IN 0 TO 30 GENERATE 
		wire_alt_sqrt_block2_w4203w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w30c_range1600w1601w4202w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w4200w(i);
	END GENERATE loop115;
	loop116 : FOR i IN 0 TO 32 GENERATE 
		wire_alt_sqrt_block2_w4280w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w32c_range1680w1681w4279w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w4277w(i);
	END GENERATE loop116;
	loop117 : FOR i IN 0 TO 34 GENERATE 
		wire_alt_sqrt_block2_w4357w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w34c_range1760w1761w4356w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w4354w(i);
	END GENERATE loop117;
	loop118 : FOR i IN 0 TO 36 GENERATE 
		wire_alt_sqrt_block2_w4434w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w36c_range1840w1841w4433w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w4431w(i);
	END GENERATE loop118;
	loop119 : FOR i IN 0 TO 38 GENERATE 
		wire_alt_sqrt_block2_w4511w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w38c_range1920w1921w4510w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w4508w(i);
	END GENERATE loop119;
	loop120 : FOR i IN 0 TO 40 GENERATE 
		wire_alt_sqrt_block2_w4588w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w40c_range2000w2001w4587w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w4585w(i);
	END GENERATE loop120;
	loop121 : FOR i IN 0 TO 42 GENERATE 
		wire_alt_sqrt_block2_w4665w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w42c_range2080w2081w4664w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w4662w(i);
	END GENERATE loop121;
	loop122 : FOR i IN 0 TO 44 GENERATE 
		wire_alt_sqrt_block2_w4742w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w44c_range2160w2161w4741w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w4739w(i);
	END GENERATE loop122;
	loop123 : FOR i IN 0 TO 46 GENERATE 
		wire_alt_sqrt_block2_w4819w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w46c_range2240w2241w4818w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w4816w(i);
	END GENERATE loop123;
	loop124 : FOR i IN 0 TO 48 GENERATE 
		wire_alt_sqrt_block2_w4896w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w48c_range2320w2321w4895w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w4893w(i);
	END GENERATE loop124;
	loop125 : FOR i IN 0 TO 5 GENERATE 
		wire_alt_sqrt_block2_w3374w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w4c_range537w538w3373w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w3371w(i);
	END GENERATE loop125;
	loop126 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w4973w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w50c_range2400w2401w4972w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w4970w(i);
	END GENERATE loop126;
	loop127 : FOR i IN 0 TO 50 GENERATE 
		wire_alt_sqrt_block2_w5051w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w52c_range448w449w5050w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w5048w(i);
	END GENERATE loop127;
	loop128 : FOR i IN 0 TO 7 GENERATE 
		wire_alt_sqrt_block2_w3436w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w6c_range619w620w3435w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w3433w(i);
	END GENERATE loop128;
	loop129 : FOR i IN 0 TO 9 GENERATE 
		wire_alt_sqrt_block2_w3498w(i) <= wire_alt_sqrt_block2_w_lg_w_lg_w_addnode_w8c_range701w702w3497w(i) OR wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w3495w(i);
	END GENERATE loop129;
	addnode_w0c <= ( wire_add_sub4_result(2 DOWNTO 0) & slevel_w0c(52 DOWNTO 0));
	addnode_w10c <= ( wire_add_sub14_result(12 DOWNTO 0) & slevel_w10c(42 DOWNTO 0));
	addnode_w11c <= ( wire_add_sub15_result(13 DOWNTO 0) & slevel_w11c(41 DOWNTO 0));
	addnode_w12c <= ( wire_add_sub16_result(14 DOWNTO 0) & slevel_w12c(40 DOWNTO 0));
	addnode_w13c <= ( wire_add_sub17_result(15 DOWNTO 0) & slevel_w13c(39 DOWNTO 0));
	addnode_w14c <= ( wire_add_sub18_result(16 DOWNTO 0) & slevel_w14c(38 DOWNTO 0));
	addnode_w15c <= ( wire_add_sub19_result(17 DOWNTO 0) & slevel_w15c(37 DOWNTO 0));
	addnode_w16c <= ( wire_add_sub20_result(18 DOWNTO 0) & slevel_w16c(36 DOWNTO 0));
	addnode_w17c <= ( wire_add_sub21_result(19 DOWNTO 0) & slevel_w17c(35 DOWNTO 0));
	addnode_w18c <= ( wire_add_sub22_result(20 DOWNTO 0) & slevel_w18c(34 DOWNTO 0));
	addnode_w19c <= ( wire_add_sub23_result(21 DOWNTO 0) & slevel_w19c(33 DOWNTO 0));
	addnode_w1c <= ( wire_add_sub5_result(3 DOWNTO 0) & slevel_w1c(51 DOWNTO 0));
	addnode_w20c <= ( wire_add_sub24_result(22 DOWNTO 0) & slevel_w20c(32 DOWNTO 0));
	addnode_w21c <= ( wire_add_sub25_result(23 DOWNTO 0) & slevel_w21c(31 DOWNTO 0));
	addnode_w22c <= ( wire_add_sub26_result(24 DOWNTO 0) & slevel_w22c(30 DOWNTO 0));
	addnode_w23c <= ( wire_add_sub27_result(25 DOWNTO 0) & slevel_w23c(29 DOWNTO 0));
	addnode_w24c <= ( wire_add_sub28_result(26 DOWNTO 0) & slevel_w24c(28 DOWNTO 0));
	addnode_w25c <= ( wire_add_sub29_result(27 DOWNTO 0) & slevel_w25c(27 DOWNTO 0));
	addnode_w26c <= ( wire_add_sub30_result(28 DOWNTO 0) & slevel_w26c(26 DOWNTO 0));
	addnode_w27c <= ( wire_add_sub31_result(27 DOWNTO 0) & qlevel_w27c(1 DOWNTO 0) & slevel_w27c(25 DOWNTO 0));
	addnode_w28c <= ( wire_add_sub32_result(27 DOWNTO 0) & "1" & qlevel_w28c(1 DOWNTO 0) & slevel_w28c(24 DOWNTO 0));
	addnode_w29c <= ( wire_add_sub33_result(28 DOWNTO 0) & "1" & qlevel_w29c(1 DOWNTO 0) & slevel_w29c(23 DOWNTO 0));
	addnode_w2c <= ( wire_add_sub6_result(4 DOWNTO 0) & slevel_w2c(50 DOWNTO 0));
	addnode_w30c <= ( wire_add_sub34_result(29 DOWNTO 0) & "1" & qlevel_w30c(1 DOWNTO 0) & slevel_w30c(22 DOWNTO 0));
	addnode_w31c <= ( wire_add_sub35_result(30 DOWNTO 0) & "1" & qlevel_w31c(1 DOWNTO 0) & slevel_w31c(21 DOWNTO 0));
	addnode_w32c <= ( wire_add_sub36_result(31 DOWNTO 0) & "1" & qlevel_w32c(1 DOWNTO 0) & slevel_w32c(20 DOWNTO 0));
	addnode_w33c <= ( wire_add_sub37_result(32 DOWNTO 0) & "1" & qlevel_w33c(1 DOWNTO 0) & slevel_w33c(19 DOWNTO 0));
	addnode_w34c <= ( wire_add_sub38_result(33 DOWNTO 0) & "1" & qlevel_w34c(1 DOWNTO 0) & slevel_w34c(18 DOWNTO 0));
	addnode_w35c <= ( wire_add_sub39_result(34 DOWNTO 0) & "1" & qlevel_w35c(1 DOWNTO 0) & slevel_w35c(17 DOWNTO 0));
	addnode_w36c <= ( wire_add_sub40_result(35 DOWNTO 0) & "1" & qlevel_w36c(1 DOWNTO 0) & slevel_w36c(16 DOWNTO 0));
	addnode_w37c <= ( wire_add_sub41_result(36 DOWNTO 0) & "1" & qlevel_w37c(1 DOWNTO 0) & slevel_w37c(15 DOWNTO 0));
	addnode_w38c <= ( wire_add_sub42_result(37 DOWNTO 0) & "1" & qlevel_w38c(1 DOWNTO 0) & slevel_w38c(14 DOWNTO 0));
	addnode_w39c <= ( wire_add_sub43_result(38 DOWNTO 0) & "1" & qlevel_w39c(1 DOWNTO 0) & slevel_w39c(13 DOWNTO 0));
	addnode_w3c <= ( wire_add_sub7_result(5 DOWNTO 0) & slevel_w3c(49 DOWNTO 0));
	addnode_w40c <= ( wire_add_sub44_result(39 DOWNTO 0) & "1" & qlevel_w40c(1 DOWNTO 0) & slevel_w40c(12 DOWNTO 0));
	addnode_w41c <= ( wire_add_sub45_result(40 DOWNTO 0) & "1" & qlevel_w41c(1 DOWNTO 0) & slevel_w41c(11 DOWNTO 0));
	addnode_w42c <= ( wire_add_sub46_result(41 DOWNTO 0) & "1" & qlevel_w42c(1 DOWNTO 0) & slevel_w42c(10 DOWNTO 0));
	addnode_w43c <= ( wire_add_sub47_result(42 DOWNTO 0) & "1" & qlevel_w43c(1 DOWNTO 0) & slevel_w43c(9 DOWNTO 0));
	addnode_w44c <= ( wire_add_sub48_result(43 DOWNTO 0) & "1" & qlevel_w44c(1 DOWNTO 0) & slevel_w44c(8 DOWNTO 0));
	addnode_w45c <= ( wire_add_sub49_result(44 DOWNTO 0) & "1" & qlevel_w45c(1 DOWNTO 0) & slevel_w45c(7 DOWNTO 0));
	addnode_w46c <= ( wire_add_sub50_result(45 DOWNTO 0) & "1" & qlevel_w46c(1 DOWNTO 0) & slevel_w46c(6 DOWNTO 0));
	addnode_w47c <= ( wire_add_sub51_result(46 DOWNTO 0) & "1" & qlevel_w47c(1 DOWNTO 0) & slevel_w47c(5 DOWNTO 0));
	addnode_w48c <= ( wire_add_sub52_result(47 DOWNTO 0) & "1" & qlevel_w48c(1 DOWNTO 0) & slevel_w48c(4 DOWNTO 0));
	addnode_w49c <= ( wire_add_sub53_result(48 DOWNTO 0) & "1" & qlevel_w49c(1 DOWNTO 0) & slevel_w49c(3 DOWNTO 0));
	addnode_w4c <= ( wire_add_sub8_result(6 DOWNTO 0) & slevel_w4c(48 DOWNTO 0));
	addnode_w50c <= ( wire_add_sub54_result(49 DOWNTO 0) & "1" & qlevel_w50c(1 DOWNTO 0) & slevel_w50c(2 DOWNTO 0));
	addnode_w51c <= ( wire_add_sub55_result(50 DOWNTO 0) & "1" & qlevel_w51c(1 DOWNTO 0) & slevel_w51c(1 DOWNTO 0));
	addnode_w52c <= ( wire_add_sub56_result(51 DOWNTO 0) & "1" & qlevel_w52c(1 DOWNTO 0) & slevel_w52c(0));
	addnode_w53c <= ( wire_add_sub57_result(52 DOWNTO 0) & "1" & qlevel_w53c(1 DOWNTO 0));
	addnode_w5c <= ( wire_add_sub9_result(7 DOWNTO 0) & slevel_w5c(47 DOWNTO 0));
	addnode_w6c <= ( wire_add_sub10_result(8 DOWNTO 0) & slevel_w6c(46 DOWNTO 0));
	addnode_w7c <= ( wire_add_sub11_result(9 DOWNTO 0) & slevel_w7c(45 DOWNTO 0));
	addnode_w8c <= ( wire_add_sub12_result(10 DOWNTO 0) & slevel_w8c(44 DOWNTO 0));
	addnode_w9c <= ( wire_add_sub13_result(11 DOWNTO 0) & slevel_w9c(43 DOWNTO 0));
	qlevel_w0c <= ( "1" & "1" & "1");
	qlevel_w10c <= ( "0" & "1" & q_ff52c(4) & q_ff50c(7 DOWNTO 6) & q_ff48c(5 DOWNTO 4) & q_ff46c(3 DOWNTO 2) & q_ff44c(1 DOWNTO 0) & "1" & "1");
	qlevel_w11c <= ( "0" & "1" & q_ff52c(4) & q_ff50c(7 DOWNTO 6) & q_ff48c(5 DOWNTO 4) & q_ff46c(3 DOWNTO 2) & q_ff44c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w784w & "1" & "1");
	qlevel_w12c <= ( "0" & "1" & q_ff52c(5) & q_ff50c(9 DOWNTO 8) & q_ff48c(7 DOWNTO 6) & q_ff46c(5 DOWNTO 4) & q_ff44c(3 DOWNTO 2) & q_ff42c(1 DOWNTO 0) & "1" & "1");
	qlevel_w13c <= ( "0" & "1" & q_ff52c(5) & q_ff50c(9 DOWNTO 8) & q_ff48c(7 DOWNTO 6) & q_ff46c(5 DOWNTO 4) & q_ff44c(3 DOWNTO 2) & q_ff42c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w866w & "1" & "1");
	qlevel_w14c <= ( "0" & "1" & q_ff52c(6) & q_ff50c(11 DOWNTO 10) & q_ff48c(9 DOWNTO 8) & q_ff46c(7 DOWNTO 6) & q_ff44c(5 DOWNTO 4) & q_ff42c(3 DOWNTO 2) & q_ff40c(1 DOWNTO 0) & "1" & "1");
	qlevel_w15c <= ( "0" & "1" & q_ff52c(6) & q_ff50c(11 DOWNTO 10) & q_ff48c(9 DOWNTO 8) & q_ff46c(7 DOWNTO 6) & q_ff44c(5 DOWNTO 4) & q_ff42c(3 DOWNTO 2) & q_ff40c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w948w & "1" & "1");
	qlevel_w16c <= ( "0" & "1" & q_ff52c(7) & q_ff50c(13 DOWNTO 12) & q_ff48c(11 DOWNTO 10) & q_ff46c(9 DOWNTO 8) & q_ff44c(7 DOWNTO 6) & q_ff42c(5 DOWNTO 4) & q_ff40c(3 DOWNTO 2) & q_ff38c(1 DOWNTO 0) & "1" & "1");
	qlevel_w17c <= ( "0" & "1" & q_ff52c(7) & q_ff50c(13 DOWNTO 12) & q_ff48c(11 DOWNTO 10) & q_ff46c(9 DOWNTO 8) & q_ff44c(7 DOWNTO 6) & q_ff42c(5 DOWNTO 4) & q_ff40c(3 DOWNTO 2) & q_ff38c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w1030w & "1" & "1");
	qlevel_w18c <= ( "0" & "1" & q_ff52c(8) & q_ff50c(15 DOWNTO 14) & q_ff48c(13 DOWNTO 12) & q_ff46c(11 DOWNTO 10) & q_ff44c(9 DOWNTO 8) & q_ff42c(7 DOWNTO 6) & q_ff40c(5 DOWNTO 4) & q_ff38c(3 DOWNTO 2) & q_ff36c(1 DOWNTO 0) & "1" & "1");
	qlevel_w19c <= ( "0" & "1" & q_ff52c(8) & q_ff50c(15 DOWNTO 14) & q_ff48c(13 DOWNTO 12) & q_ff46c(11 DOWNTO 10) & q_ff44c(9 DOWNTO 8) & q_ff42c(7 DOWNTO 6) & q_ff40c(5 DOWNTO 4) & q_ff38c(3 DOWNTO 2) & q_ff36c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w1112w & "1" & "1");
	qlevel_w1c <= ( "1" & "0" & "1" & "1");
	qlevel_w20c <= ( "0" & "1" & q_ff52c(9) & q_ff50c(17 DOWNTO 16) & q_ff48c(15 DOWNTO 14) & q_ff46c(13 DOWNTO 12) & q_ff44c(11 DOWNTO 10) & q_ff42c(9 DOWNTO 8) & q_ff40c(7 DOWNTO 6) & q_ff38c(5 DOWNTO 4) & q_ff36c(3 DOWNTO 2) & q_ff34c(1 DOWNTO 0) & "1" & "1");
	qlevel_w21c <= ( "0" & "1" & q_ff52c(9) & q_ff50c(17 DOWNTO 16) & q_ff48c(15 DOWNTO 14) & q_ff46c(13 DOWNTO 12) & q_ff44c(11 DOWNTO 10) & q_ff42c(9 DOWNTO 8) & q_ff40c(7 DOWNTO 6) & q_ff38c(5 DOWNTO 4) & q_ff36c(3 DOWNTO 2) & q_ff34c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w1194w & "1" & "1");
	qlevel_w22c <= ( "0" & "1" & q_ff52c(10) & q_ff50c(19 DOWNTO 18) & q_ff48c(17 DOWNTO 16) & q_ff46c(15 DOWNTO 14) & q_ff44c(13 DOWNTO 12) & q_ff42c(11 DOWNTO 10) & q_ff40c(9 DOWNTO 8) & q_ff38c(7 DOWNTO 6) & q_ff36c(5 DOWNTO 4) & q_ff34c(3 DOWNTO 2) & q_ff32c(1 DOWNTO 0) & "1" & "1");
	qlevel_w23c <= ( "0" & "1" & q_ff52c(10) & q_ff50c(19 DOWNTO 18) & q_ff48c(17 DOWNTO 16) & q_ff46c(15 DOWNTO 14) & q_ff44c(13 DOWNTO 12) & q_ff42c(11 DOWNTO 10) & q_ff40c(9 DOWNTO 8) & q_ff38c(7 DOWNTO 6) & q_ff36c(5 DOWNTO 4) & q_ff34c(3 DOWNTO 2) & q_ff32c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w1276w & "1" & "1");
	qlevel_w24c <= ( "0" & "1" & q_ff52c(11) & q_ff50c(21 DOWNTO 20) & q_ff48c(19 DOWNTO 18) & q_ff46c(17 DOWNTO 16) & q_ff44c(15 DOWNTO 14) & q_ff42c(13 DOWNTO 12) & q_ff40c(11 DOWNTO 10) & q_ff38c(9 DOWNTO 8) & q_ff36c(7 DOWNTO 6) & q_ff34c(5 DOWNTO 4) & q_ff32c(3 DOWNTO 2) & q_ff30c(1 DOWNTO 0) & "1" & "1");
	qlevel_w25c <= ( "0" & "1" & q_ff52c(11) & q_ff50c(21 DOWNTO 20) & q_ff48c(19 DOWNTO 18) & q_ff46c(17 DOWNTO 16) & q_ff44c(15 DOWNTO 14) & q_ff42c(13 DOWNTO 12) & q_ff40c(11 DOWNTO 10) & q_ff38c(9 DOWNTO 8) & q_ff36c(7 DOWNTO 6) & q_ff34c(5 DOWNTO 4) & q_ff32c(3 DOWNTO 2) & q_ff30c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w1358w & "1" & "1");
	qlevel_w26c <= ( "0" & "1" & q_ff52c(12) & q_ff50c(23 DOWNTO 22) & q_ff48c(21 DOWNTO 20) & q_ff46c(19 DOWNTO 18) & q_ff44c(17 DOWNTO 16) & q_ff42c(15 DOWNTO 14) & q_ff40c(13 DOWNTO 12) & q_ff38c(11 DOWNTO 10) & q_ff36c(9 DOWNTO 8) & q_ff34c(7 DOWNTO 6) & q_ff32c(5 DOWNTO 4) & q_ff30c(3 DOWNTO 2) & q_ff28c(1 DOWNTO 0) & "1" & "1");
	qlevel_w27c <= ( "0" & "1" & q_ff52c(12) & q_ff50c(23 DOWNTO 22) & q_ff48c(21 DOWNTO 20) & q_ff46c(19 DOWNTO 18) & q_ff44c(17 DOWNTO 16) & q_ff42c(15 DOWNTO 14) & q_ff40c(13 DOWNTO 12) & q_ff38c(11 DOWNTO 10) & q_ff36c(9 DOWNTO 8) & q_ff34c(7 DOWNTO 6) & q_ff32c(5 DOWNTO 4) & q_ff30c(3 DOWNTO 2) & q_ff28c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w1440w & "1" & "1");
	qlevel_w28c <= ( "0" & "1" & q_ff52c(13) & q_ff50c(25 DOWNTO 24) & q_ff48c(23 DOWNTO 22) & q_ff46c(21 DOWNTO 20) & q_ff44c(19 DOWNTO 18) & q_ff42c(17 DOWNTO 16) & q_ff40c(15 DOWNTO 14) & q_ff38c(13 DOWNTO 12) & q_ff36c(11 DOWNTO 10) & q_ff34c(9 DOWNTO 8) & q_ff32c(7 DOWNTO 6) & q_ff30c(5 DOWNTO 4) & q_ff28c(3 DOWNTO 2) & q_ff26c(1 DOWNTO 0) & "1" & "1");
	qlevel_w29c <= ( "0" & "1" & q_ff52c(13) & q_ff50c(25 DOWNTO 24) & q_ff48c(23 DOWNTO 22) & q_ff46c(21 DOWNTO 20) & q_ff44c(19 DOWNTO 18) & q_ff42c(17 DOWNTO 16) & q_ff40c(15 DOWNTO 14) & q_ff38c(13 DOWNTO 12) & q_ff36c(11 DOWNTO 10) & q_ff34c(9 DOWNTO 8) & q_ff32c(7 DOWNTO 6) & q_ff30c(5 DOWNTO 4) & q_ff28c(3 DOWNTO 2) & q_ff26c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w1521w & "1" & "1");
	qlevel_w2c <= ( "0" & "1" & q_ff52c(0) & "1" & "1");
	qlevel_w30c <= ( "0" & "1" & q_ff52c(14) & q_ff50c(27 DOWNTO 26) & q_ff48c(25 DOWNTO 24) & q_ff46c(23 DOWNTO 22) & q_ff44c(21 DOWNTO 20) & q_ff42c(19 DOWNTO 18) & q_ff40c(17 DOWNTO 16) & q_ff38c(15 DOWNTO 14) & q_ff36c(13 DOWNTO 12) & q_ff34c(11 DOWNTO 10) & q_ff32c(9 DOWNTO 8) & q_ff30c(7 DOWNTO 6) & q_ff28c(5 DOWNTO 4) & q_ff26c(3 DOWNTO 2) & q_ff24c(1 DOWNTO 0) & "1" & "1");
	qlevel_w31c <= ( "0" & "1" & q_ff52c(14) & q_ff50c(27 DOWNTO 26) & q_ff48c(25 DOWNTO 24) & q_ff46c(23 DOWNTO 22) & q_ff44c(21 DOWNTO 20) & q_ff42c(19 DOWNTO 18) & q_ff40c(17 DOWNTO 16) & q_ff38c(15 DOWNTO 14) & q_ff36c(13 DOWNTO 12) & q_ff34c(11 DOWNTO 10) & q_ff32c(9 DOWNTO 8) & q_ff30c(7 DOWNTO 6) & q_ff28c(5 DOWNTO 4) & q_ff26c(3 DOWNTO 2) & q_ff24c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w1601w & "1" & "1");
	qlevel_w32c <= ( "0" & "1" & q_ff52c(15) & q_ff50c(29 DOWNTO 28) & q_ff48c(27 DOWNTO 26) & q_ff46c(25 DOWNTO 24) & q_ff44c(23 DOWNTO 22) & q_ff42c(21 DOWNTO 20) & q_ff40c(19 DOWNTO 18) & q_ff38c(17 DOWNTO 16) & q_ff36c(15 DOWNTO 14) & q_ff34c(13 DOWNTO 12) & q_ff32c(11 DOWNTO 10) & q_ff30c(9 DOWNTO 8) & q_ff28c(7 DOWNTO 6) & q_ff26c(5 DOWNTO 4) & q_ff24c(3 DOWNTO 2) & q_ff22c(1 DOWNTO 0) & "1" & "1");
	qlevel_w33c <= ( "0" & "1" & q_ff52c(15) & q_ff50c(29 DOWNTO 28) & q_ff48c(27 DOWNTO 26) & q_ff46c(25 DOWNTO 24) & q_ff44c(23 DOWNTO 22) & q_ff42c(21 DOWNTO 20) & q_ff40c(19 DOWNTO 18) & q_ff38c(17 DOWNTO 16) & q_ff36c(15 DOWNTO 14) & q_ff34c(13 DOWNTO 12) & q_ff32c(11 DOWNTO 10) & q_ff30c(9 DOWNTO 8) & q_ff28c(7 DOWNTO 6) & q_ff26c(5 DOWNTO 4) & q_ff24c(3 DOWNTO 2) & q_ff22c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w1681w & "1" & "1");
	qlevel_w34c <= ( "0" & "1" & q_ff52c(16) & q_ff50c(31 DOWNTO 30) & q_ff48c(29 DOWNTO 28) & q_ff46c(27 DOWNTO 26) & q_ff44c(25 DOWNTO 24) & q_ff42c(23 DOWNTO 22) & q_ff40c(21 DOWNTO 20) & q_ff38c(19 DOWNTO 18) & q_ff36c(17 DOWNTO 16) & q_ff34c(15 DOWNTO 14) & q_ff32c(13 DOWNTO 12) & q_ff30c(11 DOWNTO 10) & q_ff28c(9 DOWNTO 8) & q_ff26c(7 DOWNTO 6) & q_ff24c(5 DOWNTO 4) & q_ff22c(3 DOWNTO 2) & q_ff20c(1 DOWNTO 0) & "1" & "1");
	qlevel_w35c <= ( "0" & "1" & q_ff52c(16) & q_ff50c(31 DOWNTO 30) & q_ff48c(29 DOWNTO 28) & q_ff46c(27 DOWNTO 26) & q_ff44c(25 DOWNTO 24) & q_ff42c(23 DOWNTO 22) & q_ff40c(21 DOWNTO 20) & q_ff38c(19 DOWNTO 18) & q_ff36c(17 DOWNTO 16) & q_ff34c(15 DOWNTO 14) & q_ff32c(13 DOWNTO 12) & q_ff30c(11 DOWNTO 10) & q_ff28c(9 DOWNTO 8) & q_ff26c(7 DOWNTO 6) & q_ff24c(5 DOWNTO 4) & q_ff22c(3 DOWNTO 2) & q_ff20c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w1761w & "1" & "1");
	qlevel_w36c <= ( "0" & "1" & q_ff52c(17) & q_ff50c(33 DOWNTO 32) & q_ff48c(31 DOWNTO 30) & q_ff46c(29 DOWNTO 28) & q_ff44c(27 DOWNTO 26) & q_ff42c(25 DOWNTO 24) & q_ff40c(23 DOWNTO 22) & q_ff38c(21 DOWNTO 20) & q_ff36c(19 DOWNTO 18) & q_ff34c(17 DOWNTO 16) & q_ff32c(15 DOWNTO 14) & q_ff30c(13 DOWNTO 12) & q_ff28c(11 DOWNTO 10) & q_ff26c(9 DOWNTO 8) & q_ff24c(7 DOWNTO 6) & q_ff22c(5 DOWNTO 4) & q_ff20c(3 DOWNTO 2) & q_ff18c(1 DOWNTO 0) & "1" & "1");
	qlevel_w37c <= ( "0" & "1" & q_ff52c(17) & q_ff50c(33 DOWNTO 32) & q_ff48c(31 DOWNTO 30) & q_ff46c(29 DOWNTO 28) & q_ff44c(27 DOWNTO 26) & q_ff42c(25 DOWNTO 24) & q_ff40c(23 DOWNTO 22) & q_ff38c(21 DOWNTO 20) & q_ff36c(19 DOWNTO 18) & q_ff34c(17 DOWNTO 16) & q_ff32c(15 DOWNTO 14) & q_ff30c(13 DOWNTO 12) & q_ff28c(11 DOWNTO 10) & q_ff26c(9 DOWNTO 8) & q_ff24c(7 DOWNTO 6) & q_ff22c(5 DOWNTO 4) & q_ff20c(3 DOWNTO 2) & q_ff18c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w1841w & "1" & "1");
	qlevel_w38c <= ( "0" & "1" & q_ff52c(18) & q_ff50c(35 DOWNTO 34) & q_ff48c(33 DOWNTO 32) & q_ff46c(31 DOWNTO 30) & q_ff44c(29 DOWNTO 28) & q_ff42c(27 DOWNTO 26) & q_ff40c(25 DOWNTO 24) & q_ff38c(23 DOWNTO 22) & q_ff36c(21 DOWNTO 20) & q_ff34c(19 DOWNTO 18) & q_ff32c(17 DOWNTO 16) & q_ff30c(15 DOWNTO 14) & q_ff28c(13 DOWNTO 12) & q_ff26c(11 DOWNTO 10) & q_ff24c(9 DOWNTO 8) & q_ff22c(7 DOWNTO 6) & q_ff20c(5 DOWNTO 4) & q_ff18c(3 DOWNTO 2) & q_ff16c(1 DOWNTO 0) & "1" & "1");
	qlevel_w39c <= ( "0" & "1" & q_ff52c(18) & q_ff50c(35 DOWNTO 34) & q_ff48c(33 DOWNTO 32) & q_ff46c(31 DOWNTO 30) & q_ff44c(29 DOWNTO 28) & q_ff42c(27 DOWNTO 26) & q_ff40c(25 DOWNTO 24) & q_ff38c(23 DOWNTO 22) & q_ff36c(21 DOWNTO 20) & q_ff34c(19 DOWNTO 18) & q_ff32c(17 DOWNTO 16) & q_ff30c(15 DOWNTO 14) & q_ff28c(13 DOWNTO 12) & q_ff26c(11 DOWNTO 10) & q_ff24c(9 DOWNTO 8) & q_ff22c(7 DOWNTO 6) & q_ff20c(5 DOWNTO 4) & q_ff18c(3 DOWNTO 2) & q_ff16c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w1921w & "1" & "1");
	qlevel_w3c <= ( "0" & "1" & q_ff52c(0) & wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w456w & "1" & "1");
	qlevel_w40c <= ( "0" & "1" & q_ff52c(19) & q_ff50c(37 DOWNTO 36) & q_ff48c(35 DOWNTO 34) & q_ff46c(33 DOWNTO 32) & q_ff44c(31 DOWNTO 30) & q_ff42c(29 DOWNTO 28) & q_ff40c(27 DOWNTO 26) & q_ff38c(25 DOWNTO 24) & q_ff36c(23 DOWNTO 22) & q_ff34c(21 DOWNTO 20) & q_ff32c(19 DOWNTO 18) & q_ff30c(17 DOWNTO 16) & q_ff28c(15 DOWNTO 14) & q_ff26c(13 DOWNTO 12) & q_ff24c(11 DOWNTO 10) & q_ff22c(9 DOWNTO 8) & q_ff20c(7 DOWNTO 6) & q_ff18c(5 DOWNTO 4) & q_ff16c(3 DOWNTO 2) & q_ff14c(1 DOWNTO 0) & "1" & "1");
	qlevel_w41c <= ( "0" & "1" & q_ff52c(19) & q_ff50c(37 DOWNTO 36) & q_ff48c(35 DOWNTO 34) & q_ff46c(33 DOWNTO 32) & q_ff44c(31 DOWNTO 30) & q_ff42c(29 DOWNTO 28) & q_ff40c(27 DOWNTO 26) & q_ff38c(25 DOWNTO 24) & q_ff36c(23 DOWNTO 22) & q_ff34c(21 DOWNTO 20) & q_ff32c(19 DOWNTO 18) & q_ff30c(17 DOWNTO 16) & q_ff28c(15 DOWNTO 14) & q_ff26c(13 DOWNTO 12) & q_ff24c(11 DOWNTO 10) & q_ff22c(9 DOWNTO 8) & q_ff20c(7 DOWNTO 6) & q_ff18c(5 DOWNTO 4) & q_ff16c(3 DOWNTO 2) & q_ff14c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w2001w & "1" & "1");
	qlevel_w42c <= ( "0" & "1" & q_ff52c(20) & q_ff50c(39 DOWNTO 38) & q_ff48c(37 DOWNTO 36) & q_ff46c(35 DOWNTO 34) & q_ff44c(33 DOWNTO 32) & q_ff42c(31 DOWNTO 30) & q_ff40c(29 DOWNTO 28) & q_ff38c(27 DOWNTO 26) & q_ff36c(25 DOWNTO 24) & q_ff34c(23 DOWNTO 22) & q_ff32c(21 DOWNTO 20) & q_ff30c(19 DOWNTO 18) & q_ff28c(17 DOWNTO 16) & q_ff26c(15 DOWNTO 14) & q_ff24c(13 DOWNTO 12) & q_ff22c(11 DOWNTO 10) & q_ff20c(9 DOWNTO 8) & q_ff18c(7 DOWNTO 6) & q_ff16c(5 DOWNTO 4) & q_ff14c(3 DOWNTO 2) & q_ff12c(1 DOWNTO 0) & "1" & "1");
	qlevel_w43c <= ( "0" & "1" & q_ff52c(20) & q_ff50c(39 DOWNTO 38) & q_ff48c(37 DOWNTO 36) & q_ff46c(35 DOWNTO 34) & q_ff44c(33 DOWNTO 32) & q_ff42c(31 DOWNTO 30) & q_ff40c(29 DOWNTO 28) & q_ff38c(27 DOWNTO 26) & q_ff36c(25 DOWNTO 24) & q_ff34c(23 DOWNTO 22) & q_ff32c(21 DOWNTO 20) & q_ff30c(19 DOWNTO 18) & q_ff28c(17 DOWNTO 16) & q_ff26c(15 DOWNTO 14) & q_ff24c(13 DOWNTO 12) & q_ff22c(11 DOWNTO 10) & q_ff20c(9 DOWNTO 8) & q_ff18c(7 DOWNTO 6) & q_ff16c(5 DOWNTO 4) & q_ff14c(3 DOWNTO 2) & q_ff12c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w2081w & "1" & "1");
	qlevel_w44c <= ( "0" & "1" & q_ff52c(21) & q_ff50c(41 DOWNTO 40) & q_ff48c(39 DOWNTO 38) & q_ff46c(37 DOWNTO 36) & q_ff44c(35 DOWNTO 34) & q_ff42c(33 DOWNTO 32) & q_ff40c(31 DOWNTO 30) & q_ff38c(29 DOWNTO 28) & q_ff36c(27 DOWNTO 26) & q_ff34c(25 DOWNTO 24) & q_ff32c(23 DOWNTO 22) & q_ff30c(21 DOWNTO 20) & q_ff28c(19 DOWNTO 18) & q_ff26c(17 DOWNTO 16) & q_ff24c(15 DOWNTO 14) & q_ff22c(13 DOWNTO 12) & q_ff20c(11 DOWNTO 10) & q_ff18c(9 DOWNTO 8) & q_ff16c(7 DOWNTO 6) & q_ff14c(5 DOWNTO 4) & q_ff12c(3 DOWNTO 2) & q_ff10c(1 DOWNTO 0) & "1" & "1");
	qlevel_w45c <= ( "0" & "1" & q_ff52c(21) & q_ff50c(41 DOWNTO 40) & q_ff48c(39 DOWNTO 38) & q_ff46c(37 DOWNTO 36) & q_ff44c(35 DOWNTO 34) & q_ff42c(33 DOWNTO 32) & q_ff40c(31 DOWNTO 30) & q_ff38c(29 DOWNTO 28) & q_ff36c(27 DOWNTO 26) & q_ff34c(25 DOWNTO 24) & q_ff32c(23 DOWNTO 22) & q_ff30c(21 DOWNTO 20) & q_ff28c(19 DOWNTO 18) & q_ff26c(17 DOWNTO 16) & q_ff24c(15 DOWNTO 14) & q_ff22c(13 DOWNTO 12) & q_ff20c(11 DOWNTO 10) & q_ff18c(9 DOWNTO 8) & q_ff16c(7 DOWNTO 6) & q_ff14c(5 DOWNTO 4) & q_ff12c(3 DOWNTO 2) & q_ff10c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w2161w & "1" & "1");
	qlevel_w46c <= ( "0" & "1" & q_ff52c(22) & q_ff50c(43 DOWNTO 42) & q_ff48c(41 DOWNTO 40) & q_ff46c(39 DOWNTO 38) & q_ff44c(37 DOWNTO 36) & q_ff42c(35 DOWNTO 34) & q_ff40c(33 DOWNTO 32) & q_ff38c(31 DOWNTO 30) & q_ff36c(29 DOWNTO 28) & q_ff34c(27 DOWNTO 26) & q_ff32c(25 DOWNTO 24) & q_ff30c(23 DOWNTO 22) & q_ff28c(21 DOWNTO 20) & q_ff26c(19 DOWNTO 18) & q_ff24c(17 DOWNTO 16) & q_ff22c(15 DOWNTO 14) & q_ff20c(13 DOWNTO 12) & q_ff18c(11 DOWNTO 10) & q_ff16c(9 DOWNTO 8) & q_ff14c(7 DOWNTO 6) & q_ff12c(5 DOWNTO 4) & q_ff10c(3 DOWNTO 2) & q_ff8c(1 DOWNTO 0) & "1" & "1");
	qlevel_w47c <= ( "0" & "1" & q_ff52c(22) & q_ff50c(43 DOWNTO 42) & q_ff48c(41 DOWNTO 40) & q_ff46c(39 DOWNTO 38) & q_ff44c(37 DOWNTO 36) & q_ff42c(35 DOWNTO 34) & q_ff40c(33 DOWNTO 32) & q_ff38c(31 DOWNTO 30) & q_ff36c(29 DOWNTO 28) & q_ff34c(27 DOWNTO 26) & q_ff32c(25 DOWNTO 24) & q_ff30c(23 DOWNTO 22) & q_ff28c(21 DOWNTO 20) & q_ff26c(19 DOWNTO 18) & q_ff24c(17 DOWNTO 16) & q_ff22c(15 DOWNTO 14) & q_ff20c(13 DOWNTO 12) & q_ff18c(11 DOWNTO 10) & q_ff16c(9 DOWNTO 8) & q_ff14c(7 DOWNTO 6) & q_ff12c(5 DOWNTO 4) & q_ff10c(3 DOWNTO 2) & q_ff8c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w2241w & "1" & "1");
	qlevel_w48c <= ( "0" & "1" & q_ff52c(23) & q_ff50c(45 DOWNTO 44) & q_ff48c(43 DOWNTO 42) & q_ff46c(41 DOWNTO 40) & q_ff44c(39 DOWNTO 38) & q_ff42c(37 DOWNTO 36) & q_ff40c(35 DOWNTO 34) & q_ff38c(33 DOWNTO 32) & q_ff36c(31 DOWNTO 30) & q_ff34c(29 DOWNTO 28) & q_ff32c(27 DOWNTO 26) & q_ff30c(25 DOWNTO 24) & q_ff28c(23 DOWNTO 22) & q_ff26c(21 DOWNTO 20) & q_ff24c(19 DOWNTO 18) & q_ff22c(17 DOWNTO 16) & q_ff20c(15 DOWNTO 14) & q_ff18c(13 DOWNTO 12) & q_ff16c(11 DOWNTO 10) & q_ff14c(9 DOWNTO 8) & q_ff12c(7 DOWNTO 6) & q_ff10c(5 DOWNTO 4) & q_ff8c(3 DOWNTO 2) & q_ff6c(1 DOWNTO 0) & "1" & "1");
	qlevel_w49c <= ( "0" & "1" & q_ff52c(23) & q_ff50c(45 DOWNTO 44) & q_ff48c(43 DOWNTO 42) & q_ff46c(41 DOWNTO 40) & q_ff44c(39 DOWNTO 38) & q_ff42c(37 DOWNTO 36) & q_ff40c(35 DOWNTO 34) & q_ff38c(33 DOWNTO 32) & q_ff36c(31 DOWNTO 30) & q_ff34c(29 DOWNTO 28) & q_ff32c(27 DOWNTO 26) & q_ff30c(25 DOWNTO 24) & q_ff28c(23 DOWNTO 22) & q_ff26c(21 DOWNTO 20) & q_ff24c(19 DOWNTO 18) & q_ff22c(17 DOWNTO 16) & q_ff20c(15 DOWNTO 14) & q_ff18c(13 DOWNTO 12) & q_ff16c(11 DOWNTO 10) & q_ff14c(9 DOWNTO 8) & q_ff12c(7 DOWNTO 6) & q_ff10c(5 DOWNTO 4) & q_ff8c(3 DOWNTO 2) & q_ff6c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w2321w & "1" & "1");
	qlevel_w4c <= ( "0" & "1" & q_ff52c(1) & q_ff50c(1 DOWNTO 0) & "1" & "1");
	qlevel_w50c <= ( "0" & "1" & q_ff52c(24) & q_ff50c(47 DOWNTO 46) & q_ff48c(45 DOWNTO 44) & q_ff46c(43 DOWNTO 42) & q_ff44c(41 DOWNTO 40) & q_ff42c(39 DOWNTO 38) & q_ff40c(37 DOWNTO 36) & q_ff38c(35 DOWNTO 34) & q_ff36c(33 DOWNTO 32) & q_ff34c(31 DOWNTO 30) & q_ff32c(29 DOWNTO 28) & q_ff30c(27 DOWNTO 26) & q_ff28c(25 DOWNTO 24) & q_ff26c(23 DOWNTO 22) & q_ff24c(21 DOWNTO 20) & q_ff22c(19 DOWNTO 18) & q_ff20c(17 DOWNTO 16) & q_ff18c(15 DOWNTO 14) & q_ff16c(13 DOWNTO 12) & q_ff14c(11 DOWNTO 10) & q_ff12c(9 DOWNTO 8) & q_ff10c(7 DOWNTO 6) & q_ff8c(5 DOWNTO 4) & q_ff6c(3 DOWNTO 2) & q_ff4c(1 DOWNTO 0) & "1" & "1");
	qlevel_w51c <= ( "0" & "1" & q_ff52c(24) & q_ff50c(47 DOWNTO 46) & q_ff48c(45 DOWNTO 44) & q_ff46c(43 DOWNTO 42) & q_ff44c(41 DOWNTO 40) & q_ff42c(39 DOWNTO 38) & q_ff40c(37 DOWNTO 36) & q_ff38c(35 DOWNTO 34) & q_ff36c(33 DOWNTO 32) & q_ff34c(31 DOWNTO 30) & q_ff32c(29 DOWNTO 28) & q_ff30c(27 DOWNTO 26) & q_ff28c(25 DOWNTO 24) & q_ff26c(23 DOWNTO 22) & q_ff24c(21 DOWNTO 20) & q_ff22c(19 DOWNTO 18) & q_ff20c(17 DOWNTO 16) & q_ff18c(15 DOWNTO 14) & q_ff16c(13 DOWNTO 12) & q_ff14c(11 DOWNTO 10) & q_ff12c(9 DOWNTO 8) & q_ff10c(7 DOWNTO 6) & q_ff8c(5 DOWNTO 4) & q_ff6c(3 DOWNTO 2) & q_ff4c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w2401w & "1" & "1");
	qlevel_w52c <= ( "0" & "1" & q_ff52c(25) & q_ff50c(49 DOWNTO 48) & q_ff48c(47 DOWNTO 46) & q_ff46c(45 DOWNTO 44) & q_ff44c(43 DOWNTO 42) & q_ff42c(41 DOWNTO 40) & q_ff40c(39 DOWNTO 38) & q_ff38c(37 DOWNTO 36) & q_ff36c(35 DOWNTO 34) & q_ff34c(33 DOWNTO 32) & q_ff32c(31 DOWNTO 30) & q_ff30c(29 DOWNTO 28) & q_ff28c(27 DOWNTO 26) & q_ff26c(25 DOWNTO 24) & q_ff24c(23 DOWNTO 22) & q_ff22c(21 DOWNTO 20) & q_ff20c(19 DOWNTO 18) & q_ff18c(17 DOWNTO 16) & q_ff16c(15 DOWNTO 14) & q_ff14c(13 DOWNTO 12) & q_ff12c(11 DOWNTO 10) & q_ff10c(9 DOWNTO 8) & q_ff8c(7 DOWNTO 6) & q_ff6c(5 DOWNTO 4) & q_ff4c(3 DOWNTO 2) & q_ff2c(1 DOWNTO 0) & "1" & "1");
	qlevel_w53c <= ( wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w449w & addnode_w52c(55) & q_ff52c(25) & q_ff50c(49 DOWNTO 48) & q_ff48c(47 DOWNTO 46) & q_ff46c(45 DOWNTO 44) & q_ff44c(43 DOWNTO 42) & q_ff42c(41 DOWNTO 40) & q_ff40c(39 DOWNTO 38) & q_ff38c(37 DOWNTO 36) & q_ff36c(35 DOWNTO 34) & q_ff34c(33 DOWNTO 32) & q_ff32c(31 DOWNTO 30) & q_ff30c(29 DOWNTO 28) & q_ff28c(27 DOWNTO 26) & q_ff26c(25 DOWNTO 24) & q_ff24c(23 DOWNTO 22) & q_ff22c(21 DOWNTO 20) & q_ff20c(19 DOWNTO 18) & q_ff18c(17 DOWNTO 16) & q_ff16c(15 DOWNTO 14) & q_ff14c(13 DOWNTO 12) & q_ff12c(11 DOWNTO 10) & q_ff10c(9 DOWNTO 8) & q_ff8c(7 DOWNTO 6) & q_ff6c(5 DOWNTO 4) & q_ff4c(3 DOWNTO 2) & q_ff2c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w449w & "1" & "1");
	qlevel_w5c <= ( "0" & "1" & q_ff52c(1) & q_ff50c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w538w & "1" & "1");
	qlevel_w6c <= ( "0" & "1" & q_ff52c(2) & q_ff50c(3 DOWNTO 2) & q_ff48c(1 DOWNTO 0) & "1" & "1");
	qlevel_w7c <= ( "0" & "1" & q_ff52c(2) & q_ff50c(3 DOWNTO 2) & q_ff48c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w620w & "1" & "1");
	qlevel_w8c <= ( "0" & "1" & q_ff52c(3) & q_ff50c(5 DOWNTO 4) & q_ff48c(3 DOWNTO 2) & q_ff46c(1 DOWNTO 0) & "1" & "1");
	qlevel_w9c <= ( "0" & "1" & q_ff52c(3) & q_ff50c(5 DOWNTO 4) & q_ff48c(3 DOWNTO 2) & q_ff46c(1 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w702w & "1" & "1");
	root_result <= ( "1" & q_ff52c(26) & q_ff50c(51 DOWNTO 50) & q_ff48c(49 DOWNTO 48) & q_ff46c(47 DOWNTO 46) & q_ff44c(45 DOWNTO 44) & q_ff42c(43 DOWNTO 42) & q_ff40c(41 DOWNTO 40) & q_ff38c(39 DOWNTO 38) & q_ff36c(37 DOWNTO 36) & q_ff34c(35 DOWNTO 34) & q_ff32c(33 DOWNTO 32) & q_ff30c(31 DOWNTO 30) & q_ff28c(29 DOWNTO 28) & q_ff26c(27 DOWNTO 26) & q_ff24c(25 DOWNTO 24) & q_ff22c(23 DOWNTO 22) & q_ff20c(21 DOWNTO 20) & q_ff18c(19 DOWNTO 18) & q_ff16c(17 DOWNTO 16) & q_ff14c(15 DOWNTO 14) & q_ff12c(13 DOWNTO 12) & q_ff10c(11 DOWNTO 10) & q_ff8c(9 DOWNTO 8) & q_ff6c(7 DOWNTO 6) & q_ff4c(5 DOWNTO 4) & q_ff2c(3 DOWNTO 2) & q_ff0c(1 DOWNTO 0));
	slevel_w0c <= ( "0" & rad);
	slevel_w10c <= ( rad_ff9c(44 DOWNTO 0) & "00000000000");
	slevel_w11c <= ( addnode_w10c(54 DOWNTO 11) & "000000000000");
	slevel_w12c <= ( rad_ff11c(42 DOWNTO 0) & "0000000000000");
	slevel_w13c <= ( addnode_w12c(54 DOWNTO 13) & "00000000000000");
	slevel_w14c <= ( rad_ff13c(40 DOWNTO 0) & "000000000000000");
	slevel_w15c <= ( addnode_w14c(54 DOWNTO 15) & "0000000000000000");
	slevel_w16c <= ( rad_ff15c(38 DOWNTO 0) & "00000000000000000");
	slevel_w17c <= ( addnode_w16c(54 DOWNTO 17) & "000000000000000000");
	slevel_w18c <= ( rad_ff17c(36 DOWNTO 0) & "0000000000000000000");
	slevel_w19c <= ( addnode_w18c(54 DOWNTO 19) & "00000000000000000000");
	slevel_w1c <= ( addnode_w0c(54 DOWNTO 1) & "0" & "0");
	slevel_w20c <= ( rad_ff19c(34 DOWNTO 0) & "000000000000000000000");
	slevel_w21c <= ( addnode_w20c(54 DOWNTO 21) & "0000000000000000000000");
	slevel_w22c <= ( rad_ff21c(32 DOWNTO 0) & "00000000000000000000000");
	slevel_w23c <= ( addnode_w22c(54 DOWNTO 23) & "000000000000000000000000");
	slevel_w24c <= ( rad_ff23c(30 DOWNTO 0) & "0000000000000000000000000");
	slevel_w25c <= ( addnode_w24c(54 DOWNTO 25) & "00000000000000000000000000");
	slevel_w26c <= ( rad_ff25c(28 DOWNTO 0) & "000000000000000000000000000");
	slevel_w27c <= ( addnode_w26c(54 DOWNTO 27) & "0000000000000000000000000000");
	slevel_w28c <= ( rad_ff27c(26 DOWNTO 0) & "1" & "1" & "000000000000000000000000000");
	slevel_w29c <= ( addnode_w28c(54 DOWNTO 28) & "1" & "1" & "1" & "00000000000000000000000000");
	slevel_w2c <= ( rad_ff1c(52 DOWNTO 0) & "000");
	slevel_w30c <= ( rad_ff29c(27 DOWNTO 0) & "1" & "1" & "1" & "0000000000000000000000000");
	slevel_w31c <= ( addnode_w30c(54 DOWNTO 26) & "1" & "1" & "1" & "000000000000000000000000");
	slevel_w32c <= ( rad_ff31c(29 DOWNTO 0) & "1" & "1" & "1" & "00000000000000000000000");
	slevel_w33c <= ( addnode_w32c(54 DOWNTO 24) & "1" & "1" & "1" & "0000000000000000000000");
	slevel_w34c <= ( rad_ff33c(31 DOWNTO 0) & "1" & "1" & "1" & "000000000000000000000");
	slevel_w35c <= ( addnode_w34c(54 DOWNTO 22) & "1" & "1" & "1" & "00000000000000000000");
	slevel_w36c <= ( rad_ff35c(33 DOWNTO 0) & "1" & "1" & "1" & "0000000000000000000");
	slevel_w37c <= ( addnode_w36c(54 DOWNTO 20) & "1" & "1" & "1" & "000000000000000000");
	slevel_w38c <= ( rad_ff37c(35 DOWNTO 0) & "1" & "1" & "1" & "00000000000000000");
	slevel_w39c <= ( addnode_w38c(54 DOWNTO 18) & "1" & "1" & "1" & "0000000000000000");
	slevel_w3c <= ( addnode_w2c(54 DOWNTO 3) & "0000");
	slevel_w40c <= ( rad_ff39c(37 DOWNTO 0) & "1" & "1" & "1" & "000000000000000");
	slevel_w41c <= ( addnode_w40c(54 DOWNTO 16) & "1" & "1" & "1" & "00000000000000");
	slevel_w42c <= ( rad_ff41c(39 DOWNTO 0) & "1" & "1" & "1" & "0000000000000");
	slevel_w43c <= ( addnode_w42c(54 DOWNTO 14) & "1" & "1" & "1" & "000000000000");
	slevel_w44c <= ( rad_ff43c(41 DOWNTO 0) & "1" & "1" & "1" & "00000000000");
	slevel_w45c <= ( addnode_w44c(54 DOWNTO 12) & "1" & "1" & "1" & "0000000000");
	slevel_w46c <= ( rad_ff45c(43 DOWNTO 0) & "1" & "1" & "1" & "000000000");
	slevel_w47c <= ( addnode_w46c(54 DOWNTO 10) & "1" & "1" & "1" & "00000000");
	slevel_w48c <= ( rad_ff47c(45 DOWNTO 0) & "1" & "1" & "1" & "0000000");
	slevel_w49c <= ( addnode_w48c(54 DOWNTO 8) & "1" & "1" & "1" & "000000");
	slevel_w4c <= ( rad_ff3c(50 DOWNTO 0) & "00000");
	slevel_w50c <= ( rad_ff49c(47 DOWNTO 0) & "1" & "1" & "1" & "00000");
	slevel_w51c <= ( addnode_w50c(54 DOWNTO 6) & "1" & "1" & "1" & "0000");
	slevel_w52c <= ( rad_ff51c(49 DOWNTO 0) & "1" & "1" & "1" & "000");
	slevel_w53c <= ( addnode_w52c(54 DOWNTO 4) & "1" & "1" & "1" & "00");
	slevel_w5c <= ( addnode_w4c(54 DOWNTO 5) & "000000");
	slevel_w6c <= ( rad_ff5c(48 DOWNTO 0) & "0000000");
	slevel_w7c <= ( addnode_w6c(54 DOWNTO 7) & "00000000");
	slevel_w8c <= ( rad_ff7c(46 DOWNTO 0) & "000000000");
	slevel_w9c <= ( addnode_w8c(54 DOWNTO 9) & "0000000000");
	wire_alt_sqrt_block2_w_addnode_w10c_range783w(0) <= addnode_w10c(55);
	wire_alt_sqrt_block2_w_addnode_w11c_range346w <= addnode_w11c(55 DOWNTO 12);
	wire_alt_sqrt_block2_w_addnode_w11c_range787w(0) <= addnode_w11c(55);
	wire_alt_sqrt_block2_w_addnode_w12c_range865w(0) <= addnode_w12c(55);
	wire_alt_sqrt_block2_w_addnode_w13c_range347w <= addnode_w13c(55 DOWNTO 14);
	wire_alt_sqrt_block2_w_addnode_w13c_range869w(0) <= addnode_w13c(55);
	wire_alt_sqrt_block2_w_addnode_w14c_range947w(0) <= addnode_w14c(55);
	wire_alt_sqrt_block2_w_addnode_w15c_range348w <= addnode_w15c(55 DOWNTO 16);
	wire_alt_sqrt_block2_w_addnode_w15c_range951w(0) <= addnode_w15c(55);
	wire_alt_sqrt_block2_w_addnode_w16c_range1029w(0) <= addnode_w16c(55);
	wire_alt_sqrt_block2_w_addnode_w17c_range349w <= addnode_w17c(55 DOWNTO 18);
	wire_alt_sqrt_block2_w_addnode_w17c_range1033w(0) <= addnode_w17c(55);
	wire_alt_sqrt_block2_w_addnode_w18c_range1111w(0) <= addnode_w18c(55);
	wire_alt_sqrt_block2_w_addnode_w19c_range350w <= addnode_w19c(55 DOWNTO 20);
	wire_alt_sqrt_block2_w_addnode_w19c_range1115w(0) <= addnode_w19c(55);
	wire_alt_sqrt_block2_w_addnode_w1c_range341w <= addnode_w1c(55 DOWNTO 2);
	wire_alt_sqrt_block2_w_addnode_w1c_range367w(0) <= addnode_w1c(55);
	wire_alt_sqrt_block2_w_addnode_w20c_range1193w(0) <= addnode_w20c(55);
	wire_alt_sqrt_block2_w_addnode_w21c_range351w <= addnode_w21c(55 DOWNTO 22);
	wire_alt_sqrt_block2_w_addnode_w21c_range1197w(0) <= addnode_w21c(55);
	wire_alt_sqrt_block2_w_addnode_w22c_range1275w(0) <= addnode_w22c(55);
	wire_alt_sqrt_block2_w_addnode_w23c_range352w <= addnode_w23c(55 DOWNTO 24);
	wire_alt_sqrt_block2_w_addnode_w23c_range1279w(0) <= addnode_w23c(55);
	wire_alt_sqrt_block2_w_addnode_w24c_range1357w(0) <= addnode_w24c(55);
	wire_alt_sqrt_block2_w_addnode_w25c_range353w <= addnode_w25c(55 DOWNTO 26);
	wire_alt_sqrt_block2_w_addnode_w25c_range1361w(0) <= addnode_w25c(55);
	wire_alt_sqrt_block2_w_addnode_w26c_range1439w(0) <= addnode_w26c(55);
	wire_alt_sqrt_block2_w_addnode_w27c_range354w <= addnode_w27c(55 DOWNTO 28);
	wire_alt_sqrt_block2_w_addnode_w27c_range1443w(0) <= addnode_w27c(55);
	wire_alt_sqrt_block2_w_addnode_w28c_range1520w(0) <= addnode_w28c(55);
	wire_alt_sqrt_block2_w_addnode_w29c_range355w <= addnode_w29c(55 DOWNTO 27);
	wire_alt_sqrt_block2_w_addnode_w29c_range1523w(0) <= addnode_w29c(55);
	wire_alt_sqrt_block2_w_addnode_w2c_range455w(0) <= addnode_w2c(55);
	wire_alt_sqrt_block2_w_addnode_w30c_range1600w(0) <= addnode_w30c(55);
	wire_alt_sqrt_block2_w_addnode_w31c_range356w <= addnode_w31c(55 DOWNTO 25);
	wire_alt_sqrt_block2_w_addnode_w31c_range1603w(0) <= addnode_w31c(55);
	wire_alt_sqrt_block2_w_addnode_w32c_range1680w(0) <= addnode_w32c(55);
	wire_alt_sqrt_block2_w_addnode_w33c_range357w <= addnode_w33c(55 DOWNTO 23);
	wire_alt_sqrt_block2_w_addnode_w33c_range1683w(0) <= addnode_w33c(55);
	wire_alt_sqrt_block2_w_addnode_w34c_range1760w(0) <= addnode_w34c(55);
	wire_alt_sqrt_block2_w_addnode_w35c_range358w <= addnode_w35c(55 DOWNTO 21);
	wire_alt_sqrt_block2_w_addnode_w35c_range1763w(0) <= addnode_w35c(55);
	wire_alt_sqrt_block2_w_addnode_w36c_range1840w(0) <= addnode_w36c(55);
	wire_alt_sqrt_block2_w_addnode_w37c_range359w <= addnode_w37c(55 DOWNTO 19);
	wire_alt_sqrt_block2_w_addnode_w37c_range1843w(0) <= addnode_w37c(55);
	wire_alt_sqrt_block2_w_addnode_w38c_range1920w(0) <= addnode_w38c(55);
	wire_alt_sqrt_block2_w_addnode_w39c_range360w <= addnode_w39c(55 DOWNTO 17);
	wire_alt_sqrt_block2_w_addnode_w39c_range1923w(0) <= addnode_w39c(55);
	wire_alt_sqrt_block2_w_addnode_w3c_range342w <= addnode_w3c(55 DOWNTO 4);
	wire_alt_sqrt_block2_w_addnode_w3c_range459w(0) <= addnode_w3c(55);
	wire_alt_sqrt_block2_w_addnode_w40c_range2000w(0) <= addnode_w40c(55);
	wire_alt_sqrt_block2_w_addnode_w41c_range361w <= addnode_w41c(55 DOWNTO 15);
	wire_alt_sqrt_block2_w_addnode_w41c_range2003w(0) <= addnode_w41c(55);
	wire_alt_sqrt_block2_w_addnode_w42c_range2080w(0) <= addnode_w42c(55);
	wire_alt_sqrt_block2_w_addnode_w43c_range362w <= addnode_w43c(55 DOWNTO 13);
	wire_alt_sqrt_block2_w_addnode_w43c_range2083w(0) <= addnode_w43c(55);
	wire_alt_sqrt_block2_w_addnode_w44c_range2160w(0) <= addnode_w44c(55);
	wire_alt_sqrt_block2_w_addnode_w45c_range363w <= addnode_w45c(55 DOWNTO 11);
	wire_alt_sqrt_block2_w_addnode_w45c_range2163w(0) <= addnode_w45c(55);
	wire_alt_sqrt_block2_w_addnode_w46c_range2240w(0) <= addnode_w46c(55);
	wire_alt_sqrt_block2_w_addnode_w47c_range2243w(0) <= addnode_w47c(55);
	wire_alt_sqrt_block2_w_addnode_w47c_range364w <= addnode_w47c(55 DOWNTO 9);
	wire_alt_sqrt_block2_w_addnode_w48c_range2320w(0) <= addnode_w48c(55);
	wire_alt_sqrt_block2_w_addnode_w49c_range2323w(0) <= addnode_w49c(55);
	wire_alt_sqrt_block2_w_addnode_w49c_range365w <= addnode_w49c(55 DOWNTO 7);
	wire_alt_sqrt_block2_w_addnode_w4c_range537w(0) <= addnode_w4c(55);
	wire_alt_sqrt_block2_w_addnode_w50c_range2400w(0) <= addnode_w50c(55);
	wire_alt_sqrt_block2_w_addnode_w51c_range366w <= addnode_w51c(55 DOWNTO 5);
	wire_alt_sqrt_block2_w_addnode_w51c_range2403w(0) <= addnode_w51c(55);
	wire_alt_sqrt_block2_w_addnode_w52c_range448w(0) <= addnode_w52c(55);
	wire_alt_sqrt_block2_w_addnode_w53c_range452w(0) <= addnode_w53c(55);
	wire_alt_sqrt_block2_w_addnode_w5c_range541w(0) <= addnode_w5c(55);
	wire_alt_sqrt_block2_w_addnode_w5c_range343w <= addnode_w5c(55 DOWNTO 6);
	wire_alt_sqrt_block2_w_addnode_w6c_range619w(0) <= addnode_w6c(55);
	wire_alt_sqrt_block2_w_addnode_w7c_range623w(0) <= addnode_w7c(55);
	wire_alt_sqrt_block2_w_addnode_w7c_range344w <= addnode_w7c(55 DOWNTO 8);
	wire_alt_sqrt_block2_w_addnode_w8c_range701w(0) <= addnode_w8c(55);
	wire_alt_sqrt_block2_w_addnode_w9c_range345w <= addnode_w9c(55 DOWNTO 10);
	wire_alt_sqrt_block2_w_addnode_w9c_range705w(0) <= addnode_w9c(55);
	wire_alt_sqrt_block2_w_qlevel_w10c_range3524w <= qlevel_w10c(12 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w11c_range3556w <= qlevel_w11c(13 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w12c_range3586w <= qlevel_w12c(14 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w13c_range3618w <= qlevel_w13c(15 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w14c_range3648w <= qlevel_w14c(16 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w15c_range3680w <= qlevel_w15c(17 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w16c_range3710w <= qlevel_w16c(18 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w17c_range3742w <= qlevel_w17c(19 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w18c_range3772w <= qlevel_w18c(20 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w19c_range3804w <= qlevel_w19c(21 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w20c_range3834w <= qlevel_w20c(22 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w21c_range3866w <= qlevel_w21c(23 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w22c_range3896w <= qlevel_w22c(24 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w23c_range3928w <= qlevel_w23c(25 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w24c_range3958w <= qlevel_w24c(26 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w25c_range3990w <= qlevel_w25c(27 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w26c_range4019w <= qlevel_w26c(28 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w27c_range4049w <= qlevel_w27c(29 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w28c_range4082w <= qlevel_w28c(30 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w29c_range4122w <= qlevel_w29c(31 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w2c_range3276w <= qlevel_w2c(4 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w30c_range4159w <= qlevel_w30c(32 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w31c_range4199w <= qlevel_w31c(33 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w32c_range4236w <= qlevel_w32c(34 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w33c_range4276w <= qlevel_w33c(35 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w34c_range4313w <= qlevel_w34c(36 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w35c_range4353w <= qlevel_w35c(37 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w36c_range4390w <= qlevel_w36c(38 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w37c_range4430w <= qlevel_w37c(39 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w38c_range4467w <= qlevel_w38c(40 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w39c_range4507w <= qlevel_w39c(41 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w3c_range3308w <= qlevel_w3c(5 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w40c_range4544w <= qlevel_w40c(42 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w41c_range4584w <= qlevel_w41c(43 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w42c_range4621w <= qlevel_w42c(44 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w43c_range4661w <= qlevel_w43c(45 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w44c_range4698w <= qlevel_w44c(46 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w45c_range4738w <= qlevel_w45c(47 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w46c_range4775w <= qlevel_w46c(48 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w47c_range4815w <= qlevel_w47c(49 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w48c_range4852w <= qlevel_w48c(50 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w49c_range4892w <= qlevel_w49c(51 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w4c_range3338w <= qlevel_w4c(6 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w50c_range4929w <= qlevel_w50c(52 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w51c_range4969w <= qlevel_w51c(53 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w52c_range5006w <= qlevel_w52c(54 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w53c_range5047w <= qlevel_w53c(53 DOWNTO 3);
	wire_alt_sqrt_block2_w_qlevel_w5c_range3370w <= qlevel_w5c(7 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w6c_range3400w <= qlevel_w6c(8 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w7c_range3432w <= qlevel_w7c(9 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w8c_range3462w <= qlevel_w8c(10 DOWNTO 2);
	wire_alt_sqrt_block2_w_qlevel_w9c_range3494w <= qlevel_w9c(11 DOWNTO 2);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff0c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff0c <= ( wire_alt_sqrt_block2_w_lg_w_addnode_w52c_range448w449w & wire_alt_sqrt_block2_w_lg_w_addnode_w53c_range452w453w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff10c <= ( q_ff10c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w42c_range2080w2081w & wire_alt_sqrt_block2_w_lg_w_addnode_w43c_range2083w2084w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff12c <= ( q_ff12c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w40c_range2000w2001w & wire_alt_sqrt_block2_w_lg_w_addnode_w41c_range2003w2004w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff14c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff14c <= ( q_ff14c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w38c_range1920w1921w & wire_alt_sqrt_block2_w_lg_w_addnode_w39c_range1923w1924w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff16c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff16c <= ( q_ff16c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w36c_range1840w1841w & wire_alt_sqrt_block2_w_lg_w_addnode_w37c_range1843w1844w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff18c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff18c <= ( q_ff18c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w34c_range1760w1761w & wire_alt_sqrt_block2_w_lg_w_addnode_w35c_range1763w1764w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff20c <= ( q_ff20c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w32c_range1680w1681w & wire_alt_sqrt_block2_w_lg_w_addnode_w33c_range1683w1684w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff22c <= ( q_ff22c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w30c_range1600w1601w & wire_alt_sqrt_block2_w_lg_w_addnode_w31c_range1603w1604w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff24c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff24c <= ( q_ff24c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w28c_range1520w1521w & wire_alt_sqrt_block2_w_lg_w_addnode_w29c_range1523w1524w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff26c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff26c <= ( q_ff26c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w26c_range1439w1440w & wire_alt_sqrt_block2_w_lg_w_addnode_w27c_range1443w1444w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff28c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff28c <= ( q_ff28c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w24c_range1357w1358w & wire_alt_sqrt_block2_w_lg_w_addnode_w25c_range1361w1362w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff2c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff2c <= ( q_ff2c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w50c_range2400w2401w & wire_alt_sqrt_block2_w_lg_w_addnode_w51c_range2403w2404w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff30c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff30c <= ( q_ff30c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w22c_range1275w1276w & wire_alt_sqrt_block2_w_lg_w_addnode_w23c_range1279w1280w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff32c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff32c <= ( q_ff32c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w20c_range1193w1194w & wire_alt_sqrt_block2_w_lg_w_addnode_w21c_range1197w1198w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff34c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff34c <= ( q_ff34c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w18c_range1111w1112w & wire_alt_sqrt_block2_w_lg_w_addnode_w19c_range1115w1116w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff36c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff36c <= ( q_ff36c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w16c_range1029w1030w & wire_alt_sqrt_block2_w_lg_w_addnode_w17c_range1033w1034w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff38c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff38c <= ( q_ff38c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w14c_range947w948w & wire_alt_sqrt_block2_w_lg_w_addnode_w15c_range951w952w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff40c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff40c <= ( q_ff40c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w12c_range865w866w & wire_alt_sqrt_block2_w_lg_w_addnode_w13c_range869w870w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff42c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff42c <= ( q_ff42c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w10c_range783w784w & wire_alt_sqrt_block2_w_lg_w_addnode_w11c_range787w788w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff44c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff44c <= ( q_ff44c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w8c_range701w702w & wire_alt_sqrt_block2_w_lg_w_addnode_w9c_range705w706w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff46c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff46c <= ( q_ff46c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w6c_range619w620w & wire_alt_sqrt_block2_w_lg_w_addnode_w7c_range623w624w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff48c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff48c <= ( q_ff48c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w4c_range537w538w & wire_alt_sqrt_block2_w_lg_w_addnode_w5c_range541w542w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff4c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff4c <= ( q_ff4c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w48c_range2320w2321w & wire_alt_sqrt_block2_w_lg_w_addnode_w49c_range2323w2324w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff50c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff50c <= ( q_ff50c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w2c_range455w456w & wire_alt_sqrt_block2_w_lg_w_addnode_w3c_range459w460w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff52c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff52c <= ( q_ff52c(25 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w1c_range367w368w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff6c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff6c <= ( q_ff6c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w46c_range2240w2241w & wire_alt_sqrt_block2_w_lg_w_addnode_w47c_range2243w2244w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_ff8c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_ff8c <= ( q_ff8c(49 DOWNTO 0) & wire_alt_sqrt_block2_w_lg_w_addnode_w44c_range2160w2161w & wire_alt_sqrt_block2_w_lg_w_addnode_w45c_range2163w2164w);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff11c <= wire_alt_sqrt_block2_w_addnode_w11c_range346w;
			END IF;
		END IF;
	END PROCESS;
	loop130 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff11c_w_lg_w_lg_w_q_range3587w3590w3591w(i) <= wire_rad_ff11c_w_lg_w_q_range3587w3590w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w12c_range3586w3589w(i);
	END GENERATE loop130;
	loop131 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff11c_w_lg_w_q_range3587w3588w(i) <= wire_rad_ff11c_w_q_range3587w(0) AND wire_alt_sqrt_block2_w_qlevel_w12c_range3586w(i);
	END GENERATE loop131;
	wire_rad_ff11c_w_lg_w_q_range3587w3590w(0) <= NOT wire_rad_ff11c_w_q_range3587w(0);
	loop132 : FOR i IN 0 TO 12 GENERATE 
		wire_rad_ff11c_w_lg_w_lg_w_lg_w_q_range3587w3590w3591w3592w(i) <= wire_rad_ff11c_w_lg_w_lg_w_q_range3587w3590w3591w(i) OR wire_rad_ff11c_w_lg_w_q_range3587w3588w(i);
	END GENERATE loop132;
	wire_rad_ff11c_w_q_range3587w(0) <= rad_ff11c(43);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff13c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff13c <= wire_alt_sqrt_block2_w_addnode_w13c_range347w;
			END IF;
		END IF;
	END PROCESS;
	loop133 : FOR i IN 0 TO 14 GENERATE 
		wire_rad_ff13c_w_lg_w_lg_w_q_range3649w3652w3653w(i) <= wire_rad_ff13c_w_lg_w_q_range3649w3652w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w14c_range3648w3651w(i);
	END GENERATE loop133;
	loop134 : FOR i IN 0 TO 14 GENERATE 
		wire_rad_ff13c_w_lg_w_q_range3649w3650w(i) <= wire_rad_ff13c_w_q_range3649w(0) AND wire_alt_sqrt_block2_w_qlevel_w14c_range3648w(i);
	END GENERATE loop134;
	wire_rad_ff13c_w_lg_w_q_range3649w3652w(0) <= NOT wire_rad_ff13c_w_q_range3649w(0);
	loop135 : FOR i IN 0 TO 14 GENERATE 
		wire_rad_ff13c_w_lg_w_lg_w_lg_w_q_range3649w3652w3653w3654w(i) <= wire_rad_ff13c_w_lg_w_lg_w_q_range3649w3652w3653w(i) OR wire_rad_ff13c_w_lg_w_q_range3649w3650w(i);
	END GENERATE loop135;
	wire_rad_ff13c_w_q_range3649w(0) <= rad_ff13c(41);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff15c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff15c <= wire_alt_sqrt_block2_w_addnode_w15c_range348w;
			END IF;
		END IF;
	END PROCESS;
	loop136 : FOR i IN 0 TO 16 GENERATE 
		wire_rad_ff15c_w_lg_w_lg_w_q_range3711w3714w3715w(i) <= wire_rad_ff15c_w_lg_w_q_range3711w3714w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w16c_range3710w3713w(i);
	END GENERATE loop136;
	loop137 : FOR i IN 0 TO 16 GENERATE 
		wire_rad_ff15c_w_lg_w_q_range3711w3712w(i) <= wire_rad_ff15c_w_q_range3711w(0) AND wire_alt_sqrt_block2_w_qlevel_w16c_range3710w(i);
	END GENERATE loop137;
	wire_rad_ff15c_w_lg_w_q_range3711w3714w(0) <= NOT wire_rad_ff15c_w_q_range3711w(0);
	loop138 : FOR i IN 0 TO 16 GENERATE 
		wire_rad_ff15c_w_lg_w_lg_w_lg_w_q_range3711w3714w3715w3716w(i) <= wire_rad_ff15c_w_lg_w_lg_w_q_range3711w3714w3715w(i) OR wire_rad_ff15c_w_lg_w_q_range3711w3712w(i);
	END GENERATE loop138;
	wire_rad_ff15c_w_q_range3711w(0) <= rad_ff15c(39);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff17c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff17c <= wire_alt_sqrt_block2_w_addnode_w17c_range349w;
			END IF;
		END IF;
	END PROCESS;
	loop139 : FOR i IN 0 TO 18 GENERATE 
		wire_rad_ff17c_w_lg_w_lg_w_q_range3773w3776w3777w(i) <= wire_rad_ff17c_w_lg_w_q_range3773w3776w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w18c_range3772w3775w(i);
	END GENERATE loop139;
	loop140 : FOR i IN 0 TO 18 GENERATE 
		wire_rad_ff17c_w_lg_w_q_range3773w3774w(i) <= wire_rad_ff17c_w_q_range3773w(0) AND wire_alt_sqrt_block2_w_qlevel_w18c_range3772w(i);
	END GENERATE loop140;
	wire_rad_ff17c_w_lg_w_q_range3773w3776w(0) <= NOT wire_rad_ff17c_w_q_range3773w(0);
	loop141 : FOR i IN 0 TO 18 GENERATE 
		wire_rad_ff17c_w_lg_w_lg_w_lg_w_q_range3773w3776w3777w3778w(i) <= wire_rad_ff17c_w_lg_w_lg_w_q_range3773w3776w3777w(i) OR wire_rad_ff17c_w_lg_w_q_range3773w3774w(i);
	END GENERATE loop141;
	wire_rad_ff17c_w_q_range3773w(0) <= rad_ff17c(37);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff19c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff19c <= wire_alt_sqrt_block2_w_addnode_w19c_range350w;
			END IF;
		END IF;
	END PROCESS;
	loop142 : FOR i IN 0 TO 20 GENERATE 
		wire_rad_ff19c_w_lg_w_lg_w_q_range3835w3838w3839w(i) <= wire_rad_ff19c_w_lg_w_q_range3835w3838w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w20c_range3834w3837w(i);
	END GENERATE loop142;
	loop143 : FOR i IN 0 TO 20 GENERATE 
		wire_rad_ff19c_w_lg_w_q_range3835w3836w(i) <= wire_rad_ff19c_w_q_range3835w(0) AND wire_alt_sqrt_block2_w_qlevel_w20c_range3834w(i);
	END GENERATE loop143;
	wire_rad_ff19c_w_lg_w_q_range3835w3838w(0) <= NOT wire_rad_ff19c_w_q_range3835w(0);
	loop144 : FOR i IN 0 TO 20 GENERATE 
		wire_rad_ff19c_w_lg_w_lg_w_lg_w_q_range3835w3838w3839w3840w(i) <= wire_rad_ff19c_w_lg_w_lg_w_q_range3835w3838w3839w(i) OR wire_rad_ff19c_w_lg_w_q_range3835w3836w(i);
	END GENERATE loop144;
	wire_rad_ff19c_w_q_range3835w(0) <= rad_ff19c(35);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff1c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff1c <= wire_alt_sqrt_block2_w_addnode_w1c_range341w;
			END IF;
		END IF;
	END PROCESS;
	loop145 : FOR i IN 0 TO 2 GENERATE 
		wire_rad_ff1c_w_lg_w_lg_w_q_range3277w3280w3281w(i) <= wire_rad_ff1c_w_lg_w_q_range3277w3280w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w2c_range3276w3279w(i);
	END GENERATE loop145;
	loop146 : FOR i IN 0 TO 2 GENERATE 
		wire_rad_ff1c_w_lg_w_q_range3277w3278w(i) <= wire_rad_ff1c_w_q_range3277w(0) AND wire_alt_sqrt_block2_w_qlevel_w2c_range3276w(i);
	END GENERATE loop146;
	wire_rad_ff1c_w_lg_w_q_range3277w3280w(0) <= NOT wire_rad_ff1c_w_q_range3277w(0);
	loop147 : FOR i IN 0 TO 2 GENERATE 
		wire_rad_ff1c_w_lg_w_lg_w_lg_w_q_range3277w3280w3281w3282w(i) <= wire_rad_ff1c_w_lg_w_lg_w_q_range3277w3280w3281w(i) OR wire_rad_ff1c_w_lg_w_q_range3277w3278w(i);
	END GENERATE loop147;
	wire_rad_ff1c_w_q_range3277w(0) <= rad_ff1c(53);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff21c <= wire_alt_sqrt_block2_w_addnode_w21c_range351w;
			END IF;
		END IF;
	END PROCESS;
	loop148 : FOR i IN 0 TO 22 GENERATE 
		wire_rad_ff21c_w_lg_w_lg_w_q_range3897w3900w3901w(i) <= wire_rad_ff21c_w_lg_w_q_range3897w3900w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w22c_range3896w3899w(i);
	END GENERATE loop148;
	loop149 : FOR i IN 0 TO 22 GENERATE 
		wire_rad_ff21c_w_lg_w_q_range3897w3898w(i) <= wire_rad_ff21c_w_q_range3897w(0) AND wire_alt_sqrt_block2_w_qlevel_w22c_range3896w(i);
	END GENERATE loop149;
	wire_rad_ff21c_w_lg_w_q_range3897w3900w(0) <= NOT wire_rad_ff21c_w_q_range3897w(0);
	loop150 : FOR i IN 0 TO 22 GENERATE 
		wire_rad_ff21c_w_lg_w_lg_w_lg_w_q_range3897w3900w3901w3902w(i) <= wire_rad_ff21c_w_lg_w_lg_w_q_range3897w3900w3901w(i) OR wire_rad_ff21c_w_lg_w_q_range3897w3898w(i);
	END GENERATE loop150;
	wire_rad_ff21c_w_q_range3897w(0) <= rad_ff21c(33);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff23c <= wire_alt_sqrt_block2_w_addnode_w23c_range352w;
			END IF;
		END IF;
	END PROCESS;
	loop151 : FOR i IN 0 TO 24 GENERATE 
		wire_rad_ff23c_w_lg_w_lg_w_q_range3959w3962w3963w(i) <= wire_rad_ff23c_w_lg_w_q_range3959w3962w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w24c_range3958w3961w(i);
	END GENERATE loop151;
	loop152 : FOR i IN 0 TO 24 GENERATE 
		wire_rad_ff23c_w_lg_w_q_range3959w3960w(i) <= wire_rad_ff23c_w_q_range3959w(0) AND wire_alt_sqrt_block2_w_qlevel_w24c_range3958w(i);
	END GENERATE loop152;
	wire_rad_ff23c_w_lg_w_q_range3959w3962w(0) <= NOT wire_rad_ff23c_w_q_range3959w(0);
	loop153 : FOR i IN 0 TO 24 GENERATE 
		wire_rad_ff23c_w_lg_w_lg_w_lg_w_q_range3959w3962w3963w3964w(i) <= wire_rad_ff23c_w_lg_w_lg_w_q_range3959w3962w3963w(i) OR wire_rad_ff23c_w_lg_w_q_range3959w3960w(i);
	END GENERATE loop153;
	wire_rad_ff23c_w_q_range3959w(0) <= rad_ff23c(31);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff25c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff25c <= wire_alt_sqrt_block2_w_addnode_w25c_range353w;
			END IF;
		END IF;
	END PROCESS;
	loop154 : FOR i IN 0 TO 26 GENERATE 
		wire_rad_ff25c_w_lg_w_lg_w_q_range4020w4023w4024w(i) <= wire_rad_ff25c_w_lg_w_q_range4020w4023w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w26c_range4019w4022w(i);
	END GENERATE loop154;
	loop155 : FOR i IN 0 TO 26 GENERATE 
		wire_rad_ff25c_w_lg_w_q_range4020w4021w(i) <= wire_rad_ff25c_w_q_range4020w(0) AND wire_alt_sqrt_block2_w_qlevel_w26c_range4019w(i);
	END GENERATE loop155;
	wire_rad_ff25c_w_lg_w_q_range4020w4023w(0) <= NOT wire_rad_ff25c_w_q_range4020w(0);
	loop156 : FOR i IN 0 TO 26 GENERATE 
		wire_rad_ff25c_w_lg_w_lg_w_lg_w_q_range4020w4023w4024w4025w(i) <= wire_rad_ff25c_w_lg_w_lg_w_q_range4020w4023w4024w(i) OR wire_rad_ff25c_w_lg_w_q_range4020w4021w(i);
	END GENERATE loop156;
	wire_rad_ff25c_w_q_range4020w(0) <= rad_ff25c(29);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff27c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff27c <= wire_alt_sqrt_block2_w_addnode_w27c_range354w;
			END IF;
		END IF;
	END PROCESS;
	loop157 : FOR i IN 0 TO 27 GENERATE 
		wire_rad_ff27c_w_lg_w_lg_w_q_range4083w4086w4087w(i) <= wire_rad_ff27c_w_lg_w_q_range4083w4086w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w28c_range4082w4085w(i);
	END GENERATE loop157;
	loop158 : FOR i IN 0 TO 27 GENERATE 
		wire_rad_ff27c_w_lg_w_q_range4083w4084w(i) <= wire_rad_ff27c_w_q_range4083w(0) AND wire_alt_sqrt_block2_w_qlevel_w28c_range4082w(i);
	END GENERATE loop158;
	wire_rad_ff27c_w_lg_w_q_range4083w4086w(0) <= NOT wire_rad_ff27c_w_q_range4083w(0);
	loop159 : FOR i IN 0 TO 27 GENERATE 
		wire_rad_ff27c_w_lg_w_lg_w_lg_w_q_range4083w4086w4087w4088w(i) <= wire_rad_ff27c_w_lg_w_lg_w_q_range4083w4086w4087w(i) OR wire_rad_ff27c_w_lg_w_q_range4083w4084w(i);
	END GENERATE loop159;
	wire_rad_ff27c_w_q_range4083w(0) <= rad_ff27c(27);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff29c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff29c <= wire_alt_sqrt_block2_w_addnode_w29c_range355w;
			END IF;
		END IF;
	END PROCESS;
	loop160 : FOR i IN 0 TO 29 GENERATE 
		wire_rad_ff29c_w_lg_w_lg_w_q_range4160w4163w4164w(i) <= wire_rad_ff29c_w_lg_w_q_range4160w4163w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w30c_range4159w4162w(i);
	END GENERATE loop160;
	loop161 : FOR i IN 0 TO 29 GENERATE 
		wire_rad_ff29c_w_lg_w_q_range4160w4161w(i) <= wire_rad_ff29c_w_q_range4160w(0) AND wire_alt_sqrt_block2_w_qlevel_w30c_range4159w(i);
	END GENERATE loop161;
	wire_rad_ff29c_w_lg_w_q_range4160w4163w(0) <= NOT wire_rad_ff29c_w_q_range4160w(0);
	loop162 : FOR i IN 0 TO 29 GENERATE 
		wire_rad_ff29c_w_lg_w_lg_w_lg_w_q_range4160w4163w4164w4165w(i) <= wire_rad_ff29c_w_lg_w_lg_w_q_range4160w4163w4164w(i) OR wire_rad_ff29c_w_lg_w_q_range4160w4161w(i);
	END GENERATE loop162;
	wire_rad_ff29c_w_q_range4160w(0) <= rad_ff29c(28);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff31c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff31c <= wire_alt_sqrt_block2_w_addnode_w31c_range356w;
			END IF;
		END IF;
	END PROCESS;
	loop163 : FOR i IN 0 TO 31 GENERATE 
		wire_rad_ff31c_w_lg_w_lg_w_q_range4237w4240w4241w(i) <= wire_rad_ff31c_w_lg_w_q_range4237w4240w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w32c_range4236w4239w(i);
	END GENERATE loop163;
	loop164 : FOR i IN 0 TO 31 GENERATE 
		wire_rad_ff31c_w_lg_w_q_range4237w4238w(i) <= wire_rad_ff31c_w_q_range4237w(0) AND wire_alt_sqrt_block2_w_qlevel_w32c_range4236w(i);
	END GENERATE loop164;
	wire_rad_ff31c_w_lg_w_q_range4237w4240w(0) <= NOT wire_rad_ff31c_w_q_range4237w(0);
	loop165 : FOR i IN 0 TO 31 GENERATE 
		wire_rad_ff31c_w_lg_w_lg_w_lg_w_q_range4237w4240w4241w4242w(i) <= wire_rad_ff31c_w_lg_w_lg_w_q_range4237w4240w4241w(i) OR wire_rad_ff31c_w_lg_w_q_range4237w4238w(i);
	END GENERATE loop165;
	wire_rad_ff31c_w_q_range4237w(0) <= rad_ff31c(30);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff33c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff33c <= wire_alt_sqrt_block2_w_addnode_w33c_range357w;
			END IF;
		END IF;
	END PROCESS;
	loop166 : FOR i IN 0 TO 33 GENERATE 
		wire_rad_ff33c_w_lg_w_lg_w_q_range4314w4317w4318w(i) <= wire_rad_ff33c_w_lg_w_q_range4314w4317w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w34c_range4313w4316w(i);
	END GENERATE loop166;
	loop167 : FOR i IN 0 TO 33 GENERATE 
		wire_rad_ff33c_w_lg_w_q_range4314w4315w(i) <= wire_rad_ff33c_w_q_range4314w(0) AND wire_alt_sqrt_block2_w_qlevel_w34c_range4313w(i);
	END GENERATE loop167;
	wire_rad_ff33c_w_lg_w_q_range4314w4317w(0) <= NOT wire_rad_ff33c_w_q_range4314w(0);
	loop168 : FOR i IN 0 TO 33 GENERATE 
		wire_rad_ff33c_w_lg_w_lg_w_lg_w_q_range4314w4317w4318w4319w(i) <= wire_rad_ff33c_w_lg_w_lg_w_q_range4314w4317w4318w(i) OR wire_rad_ff33c_w_lg_w_q_range4314w4315w(i);
	END GENERATE loop168;
	wire_rad_ff33c_w_q_range4314w(0) <= rad_ff33c(32);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff35c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff35c <= wire_alt_sqrt_block2_w_addnode_w35c_range358w;
			END IF;
		END IF;
	END PROCESS;
	loop169 : FOR i IN 0 TO 35 GENERATE 
		wire_rad_ff35c_w_lg_w_lg_w_q_range4391w4394w4395w(i) <= wire_rad_ff35c_w_lg_w_q_range4391w4394w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w36c_range4390w4393w(i);
	END GENERATE loop169;
	loop170 : FOR i IN 0 TO 35 GENERATE 
		wire_rad_ff35c_w_lg_w_q_range4391w4392w(i) <= wire_rad_ff35c_w_q_range4391w(0) AND wire_alt_sqrt_block2_w_qlevel_w36c_range4390w(i);
	END GENERATE loop170;
	wire_rad_ff35c_w_lg_w_q_range4391w4394w(0) <= NOT wire_rad_ff35c_w_q_range4391w(0);
	loop171 : FOR i IN 0 TO 35 GENERATE 
		wire_rad_ff35c_w_lg_w_lg_w_lg_w_q_range4391w4394w4395w4396w(i) <= wire_rad_ff35c_w_lg_w_lg_w_q_range4391w4394w4395w(i) OR wire_rad_ff35c_w_lg_w_q_range4391w4392w(i);
	END GENERATE loop171;
	wire_rad_ff35c_w_q_range4391w(0) <= rad_ff35c(34);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff37c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff37c <= wire_alt_sqrt_block2_w_addnode_w37c_range359w;
			END IF;
		END IF;
	END PROCESS;
	loop172 : FOR i IN 0 TO 37 GENERATE 
		wire_rad_ff37c_w_lg_w_lg_w_q_range4468w4471w4472w(i) <= wire_rad_ff37c_w_lg_w_q_range4468w4471w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w38c_range4467w4470w(i);
	END GENERATE loop172;
	loop173 : FOR i IN 0 TO 37 GENERATE 
		wire_rad_ff37c_w_lg_w_q_range4468w4469w(i) <= wire_rad_ff37c_w_q_range4468w(0) AND wire_alt_sqrt_block2_w_qlevel_w38c_range4467w(i);
	END GENERATE loop173;
	wire_rad_ff37c_w_lg_w_q_range4468w4471w(0) <= NOT wire_rad_ff37c_w_q_range4468w(0);
	loop174 : FOR i IN 0 TO 37 GENERATE 
		wire_rad_ff37c_w_lg_w_lg_w_lg_w_q_range4468w4471w4472w4473w(i) <= wire_rad_ff37c_w_lg_w_lg_w_q_range4468w4471w4472w(i) OR wire_rad_ff37c_w_lg_w_q_range4468w4469w(i);
	END GENERATE loop174;
	wire_rad_ff37c_w_q_range4468w(0) <= rad_ff37c(36);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff39c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff39c <= wire_alt_sqrt_block2_w_addnode_w39c_range360w;
			END IF;
		END IF;
	END PROCESS;
	loop175 : FOR i IN 0 TO 39 GENERATE 
		wire_rad_ff39c_w_lg_w_lg_w_q_range4545w4548w4549w(i) <= wire_rad_ff39c_w_lg_w_q_range4545w4548w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w40c_range4544w4547w(i);
	END GENERATE loop175;
	loop176 : FOR i IN 0 TO 39 GENERATE 
		wire_rad_ff39c_w_lg_w_q_range4545w4546w(i) <= wire_rad_ff39c_w_q_range4545w(0) AND wire_alt_sqrt_block2_w_qlevel_w40c_range4544w(i);
	END GENERATE loop176;
	wire_rad_ff39c_w_lg_w_q_range4545w4548w(0) <= NOT wire_rad_ff39c_w_q_range4545w(0);
	loop177 : FOR i IN 0 TO 39 GENERATE 
		wire_rad_ff39c_w_lg_w_lg_w_lg_w_q_range4545w4548w4549w4550w(i) <= wire_rad_ff39c_w_lg_w_lg_w_q_range4545w4548w4549w(i) OR wire_rad_ff39c_w_lg_w_q_range4545w4546w(i);
	END GENERATE loop177;
	wire_rad_ff39c_w_q_range4545w(0) <= rad_ff39c(38);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff3c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff3c <= wire_alt_sqrt_block2_w_addnode_w3c_range342w;
			END IF;
		END IF;
	END PROCESS;
	loop178 : FOR i IN 0 TO 4 GENERATE 
		wire_rad_ff3c_w_lg_w_lg_w_q_range3339w3342w3343w(i) <= wire_rad_ff3c_w_lg_w_q_range3339w3342w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w4c_range3338w3341w(i);
	END GENERATE loop178;
	loop179 : FOR i IN 0 TO 4 GENERATE 
		wire_rad_ff3c_w_lg_w_q_range3339w3340w(i) <= wire_rad_ff3c_w_q_range3339w(0) AND wire_alt_sqrt_block2_w_qlevel_w4c_range3338w(i);
	END GENERATE loop179;
	wire_rad_ff3c_w_lg_w_q_range3339w3342w(0) <= NOT wire_rad_ff3c_w_q_range3339w(0);
	loop180 : FOR i IN 0 TO 4 GENERATE 
		wire_rad_ff3c_w_lg_w_lg_w_lg_w_q_range3339w3342w3343w3344w(i) <= wire_rad_ff3c_w_lg_w_lg_w_q_range3339w3342w3343w(i) OR wire_rad_ff3c_w_lg_w_q_range3339w3340w(i);
	END GENERATE loop180;
	wire_rad_ff3c_w_q_range3339w(0) <= rad_ff3c(51);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff41c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff41c <= wire_alt_sqrt_block2_w_addnode_w41c_range361w;
			END IF;
		END IF;
	END PROCESS;
	loop181 : FOR i IN 0 TO 41 GENERATE 
		wire_rad_ff41c_w_lg_w_lg_w_q_range4622w4625w4626w(i) <= wire_rad_ff41c_w_lg_w_q_range4622w4625w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w42c_range4621w4624w(i);
	END GENERATE loop181;
	loop182 : FOR i IN 0 TO 41 GENERATE 
		wire_rad_ff41c_w_lg_w_q_range4622w4623w(i) <= wire_rad_ff41c_w_q_range4622w(0) AND wire_alt_sqrt_block2_w_qlevel_w42c_range4621w(i);
	END GENERATE loop182;
	wire_rad_ff41c_w_lg_w_q_range4622w4625w(0) <= NOT wire_rad_ff41c_w_q_range4622w(0);
	loop183 : FOR i IN 0 TO 41 GENERATE 
		wire_rad_ff41c_w_lg_w_lg_w_lg_w_q_range4622w4625w4626w4627w(i) <= wire_rad_ff41c_w_lg_w_lg_w_q_range4622w4625w4626w(i) OR wire_rad_ff41c_w_lg_w_q_range4622w4623w(i);
	END GENERATE loop183;
	wire_rad_ff41c_w_q_range4622w(0) <= rad_ff41c(40);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff43c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff43c <= wire_alt_sqrt_block2_w_addnode_w43c_range362w;
			END IF;
		END IF;
	END PROCESS;
	loop184 : FOR i IN 0 TO 43 GENERATE 
		wire_rad_ff43c_w_lg_w_lg_w_q_range4699w4702w4703w(i) <= wire_rad_ff43c_w_lg_w_q_range4699w4702w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w44c_range4698w4701w(i);
	END GENERATE loop184;
	loop185 : FOR i IN 0 TO 43 GENERATE 
		wire_rad_ff43c_w_lg_w_q_range4699w4700w(i) <= wire_rad_ff43c_w_q_range4699w(0) AND wire_alt_sqrt_block2_w_qlevel_w44c_range4698w(i);
	END GENERATE loop185;
	wire_rad_ff43c_w_lg_w_q_range4699w4702w(0) <= NOT wire_rad_ff43c_w_q_range4699w(0);
	loop186 : FOR i IN 0 TO 43 GENERATE 
		wire_rad_ff43c_w_lg_w_lg_w_lg_w_q_range4699w4702w4703w4704w(i) <= wire_rad_ff43c_w_lg_w_lg_w_q_range4699w4702w4703w(i) OR wire_rad_ff43c_w_lg_w_q_range4699w4700w(i);
	END GENERATE loop186;
	wire_rad_ff43c_w_q_range4699w(0) <= rad_ff43c(42);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff45c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff45c <= wire_alt_sqrt_block2_w_addnode_w45c_range363w;
			END IF;
		END IF;
	END PROCESS;
	loop187 : FOR i IN 0 TO 45 GENERATE 
		wire_rad_ff45c_w_lg_w_lg_w_q_range4776w4779w4780w(i) <= wire_rad_ff45c_w_lg_w_q_range4776w4779w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w46c_range4775w4778w(i);
	END GENERATE loop187;
	loop188 : FOR i IN 0 TO 45 GENERATE 
		wire_rad_ff45c_w_lg_w_q_range4776w4777w(i) <= wire_rad_ff45c_w_q_range4776w(0) AND wire_alt_sqrt_block2_w_qlevel_w46c_range4775w(i);
	END GENERATE loop188;
	wire_rad_ff45c_w_lg_w_q_range4776w4779w(0) <= NOT wire_rad_ff45c_w_q_range4776w(0);
	loop189 : FOR i IN 0 TO 45 GENERATE 
		wire_rad_ff45c_w_lg_w_lg_w_lg_w_q_range4776w4779w4780w4781w(i) <= wire_rad_ff45c_w_lg_w_lg_w_q_range4776w4779w4780w(i) OR wire_rad_ff45c_w_lg_w_q_range4776w4777w(i);
	END GENERATE loop189;
	wire_rad_ff45c_w_q_range4776w(0) <= rad_ff45c(44);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff47c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff47c <= wire_alt_sqrt_block2_w_addnode_w47c_range364w;
			END IF;
		END IF;
	END PROCESS;
	loop190 : FOR i IN 0 TO 47 GENERATE 
		wire_rad_ff47c_w_lg_w_lg_w_q_range4853w4856w4857w(i) <= wire_rad_ff47c_w_lg_w_q_range4853w4856w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w48c_range4852w4855w(i);
	END GENERATE loop190;
	loop191 : FOR i IN 0 TO 47 GENERATE 
		wire_rad_ff47c_w_lg_w_q_range4853w4854w(i) <= wire_rad_ff47c_w_q_range4853w(0) AND wire_alt_sqrt_block2_w_qlevel_w48c_range4852w(i);
	END GENERATE loop191;
	wire_rad_ff47c_w_lg_w_q_range4853w4856w(0) <= NOT wire_rad_ff47c_w_q_range4853w(0);
	loop192 : FOR i IN 0 TO 47 GENERATE 
		wire_rad_ff47c_w_lg_w_lg_w_lg_w_q_range4853w4856w4857w4858w(i) <= wire_rad_ff47c_w_lg_w_lg_w_q_range4853w4856w4857w(i) OR wire_rad_ff47c_w_lg_w_q_range4853w4854w(i);
	END GENERATE loop192;
	wire_rad_ff47c_w_q_range4853w(0) <= rad_ff47c(46);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff49c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff49c <= wire_alt_sqrt_block2_w_addnode_w49c_range365w;
			END IF;
		END IF;
	END PROCESS;
	loop193 : FOR i IN 0 TO 49 GENERATE 
		wire_rad_ff49c_w_lg_w_lg_w_q_range4930w4933w4934w(i) <= wire_rad_ff49c_w_lg_w_q_range4930w4933w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w50c_range4929w4932w(i);
	END GENERATE loop193;
	loop194 : FOR i IN 0 TO 49 GENERATE 
		wire_rad_ff49c_w_lg_w_q_range4930w4931w(i) <= wire_rad_ff49c_w_q_range4930w(0) AND wire_alt_sqrt_block2_w_qlevel_w50c_range4929w(i);
	END GENERATE loop194;
	wire_rad_ff49c_w_lg_w_q_range4930w4933w(0) <= NOT wire_rad_ff49c_w_q_range4930w(0);
	loop195 : FOR i IN 0 TO 49 GENERATE 
		wire_rad_ff49c_w_lg_w_lg_w_lg_w_q_range4930w4933w4934w4935w(i) <= wire_rad_ff49c_w_lg_w_lg_w_q_range4930w4933w4934w(i) OR wire_rad_ff49c_w_lg_w_q_range4930w4931w(i);
	END GENERATE loop195;
	wire_rad_ff49c_w_q_range4930w(0) <= rad_ff49c(48);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff51c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff51c <= wire_alt_sqrt_block2_w_addnode_w51c_range366w;
			END IF;
		END IF;
	END PROCESS;
	loop196 : FOR i IN 0 TO 51 GENERATE 
		wire_rad_ff51c_w_lg_w_lg_w_q_range5007w5010w5011w(i) <= wire_rad_ff51c_w_lg_w_q_range5007w5010w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w52c_range5006w5009w(i);
	END GENERATE loop196;
	loop197 : FOR i IN 0 TO 51 GENERATE 
		wire_rad_ff51c_w_lg_w_q_range5007w5008w(i) <= wire_rad_ff51c_w_q_range5007w(0) AND wire_alt_sqrt_block2_w_qlevel_w52c_range5006w(i);
	END GENERATE loop197;
	wire_rad_ff51c_w_lg_w_q_range5007w5010w(0) <= NOT wire_rad_ff51c_w_q_range5007w(0);
	loop198 : FOR i IN 0 TO 51 GENERATE 
		wire_rad_ff51c_w_lg_w_lg_w_lg_w_q_range5007w5010w5011w5012w(i) <= wire_rad_ff51c_w_lg_w_lg_w_q_range5007w5010w5011w(i) OR wire_rad_ff51c_w_lg_w_q_range5007w5008w(i);
	END GENERATE loop198;
	wire_rad_ff51c_w_q_range5007w(0) <= rad_ff51c(50);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff5c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff5c <= wire_alt_sqrt_block2_w_addnode_w5c_range343w;
			END IF;
		END IF;
	END PROCESS;
	loop199 : FOR i IN 0 TO 6 GENERATE 
		wire_rad_ff5c_w_lg_w_lg_w_q_range3401w3404w3405w(i) <= wire_rad_ff5c_w_lg_w_q_range3401w3404w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w6c_range3400w3403w(i);
	END GENERATE loop199;
	loop200 : FOR i IN 0 TO 6 GENERATE 
		wire_rad_ff5c_w_lg_w_q_range3401w3402w(i) <= wire_rad_ff5c_w_q_range3401w(0) AND wire_alt_sqrt_block2_w_qlevel_w6c_range3400w(i);
	END GENERATE loop200;
	wire_rad_ff5c_w_lg_w_q_range3401w3404w(0) <= NOT wire_rad_ff5c_w_q_range3401w(0);
	loop201 : FOR i IN 0 TO 6 GENERATE 
		wire_rad_ff5c_w_lg_w_lg_w_lg_w_q_range3401w3404w3405w3406w(i) <= wire_rad_ff5c_w_lg_w_lg_w_q_range3401w3404w3405w(i) OR wire_rad_ff5c_w_lg_w_q_range3401w3402w(i);
	END GENERATE loop201;
	wire_rad_ff5c_w_q_range3401w(0) <= rad_ff5c(49);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff7c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff7c <= wire_alt_sqrt_block2_w_addnode_w7c_range344w;
			END IF;
		END IF;
	END PROCESS;
	loop202 : FOR i IN 0 TO 8 GENERATE 
		wire_rad_ff7c_w_lg_w_lg_w_q_range3463w3466w3467w(i) <= wire_rad_ff7c_w_lg_w_q_range3463w3466w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w8c_range3462w3465w(i);
	END GENERATE loop202;
	loop203 : FOR i IN 0 TO 8 GENERATE 
		wire_rad_ff7c_w_lg_w_q_range3463w3464w(i) <= wire_rad_ff7c_w_q_range3463w(0) AND wire_alt_sqrt_block2_w_qlevel_w8c_range3462w(i);
	END GENERATE loop203;
	wire_rad_ff7c_w_lg_w_q_range3463w3466w(0) <= NOT wire_rad_ff7c_w_q_range3463w(0);
	loop204 : FOR i IN 0 TO 8 GENERATE 
		wire_rad_ff7c_w_lg_w_lg_w_lg_w_q_range3463w3466w3467w3468w(i) <= wire_rad_ff7c_w_lg_w_lg_w_q_range3463w3466w3467w(i) OR wire_rad_ff7c_w_lg_w_q_range3463w3464w(i);
	END GENERATE loop204;
	wire_rad_ff7c_w_q_range3463w(0) <= rad_ff7c(47);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rad_ff9c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rad_ff9c <= wire_alt_sqrt_block2_w_addnode_w9c_range345w;
			END IF;
		END IF;
	END PROCESS;
	loop205 : FOR i IN 0 TO 10 GENERATE 
		wire_rad_ff9c_w_lg_w_lg_w_q_range3525w3528w3529w(i) <= wire_rad_ff9c_w_lg_w_q_range3525w3528w(0) AND wire_alt_sqrt_block2_w_lg_w_qlevel_w10c_range3524w3527w(i);
	END GENERATE loop205;
	loop206 : FOR i IN 0 TO 10 GENERATE 
		wire_rad_ff9c_w_lg_w_q_range3525w3526w(i) <= wire_rad_ff9c_w_q_range3525w(0) AND wire_alt_sqrt_block2_w_qlevel_w10c_range3524w(i);
	END GENERATE loop206;
	wire_rad_ff9c_w_lg_w_q_range3525w3528w(0) <= NOT wire_rad_ff9c_w_q_range3525w(0);
	loop207 : FOR i IN 0 TO 10 GENERATE 
		wire_rad_ff9c_w_lg_w_lg_w_lg_w_q_range3525w3528w3529w3530w(i) <= wire_rad_ff9c_w_lg_w_lg_w_q_range3525w3528w3529w(i) OR wire_rad_ff9c_w_lg_w_q_range3525w3526w(i);
	END GENERATE loop207;
	wire_rad_ff9c_w_q_range3525w(0) <= rad_ff9c(45);
	wire_add_sub10_dataa <= ( slevel_w6c(55 DOWNTO 47));
	wire_add_sub10_datab <= ( wire_rad_ff5c_w_lg_w_lg_w_lg_w_q_range3401w3404w3405w3406w & qlevel_w6c(1 DOWNTO 0));
	add_sub10 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => wire_add_sub10_dataa,
		datab => wire_add_sub10_datab,
		result => wire_add_sub10_result
	  );
	wire_add_sub11_dataa <= ( slevel_w7c(55 DOWNTO 46));
	wire_add_sub11_datab <= ( wire_alt_sqrt_block2_w3436w & qlevel_w7c(1 DOWNTO 0));
	add_sub11 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 10
	  )
	  PORT MAP ( 
		dataa => wire_add_sub11_dataa,
		datab => wire_add_sub11_datab,
		result => wire_add_sub11_result
	  );
	wire_add_sub12_dataa <= ( slevel_w8c(55 DOWNTO 45));
	wire_add_sub12_datab <= ( wire_rad_ff7c_w_lg_w_lg_w_lg_w_q_range3463w3466w3467w3468w & qlevel_w8c(1 DOWNTO 0));
	add_sub12 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 11
	  )
	  PORT MAP ( 
		dataa => wire_add_sub12_dataa,
		datab => wire_add_sub12_datab,
		result => wire_add_sub12_result
	  );
	wire_add_sub13_dataa <= ( slevel_w9c(55 DOWNTO 44));
	wire_add_sub13_datab <= ( wire_alt_sqrt_block2_w3498w & qlevel_w9c(1 DOWNTO 0));
	add_sub13 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => wire_add_sub13_dataa,
		datab => wire_add_sub13_datab,
		result => wire_add_sub13_result
	  );
	wire_add_sub14_dataa <= ( slevel_w10c(55 DOWNTO 43));
	wire_add_sub14_datab <= ( wire_rad_ff9c_w_lg_w_lg_w_lg_w_q_range3525w3528w3529w3530w & qlevel_w10c(1 DOWNTO 0));
	add_sub14 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		dataa => wire_add_sub14_dataa,
		datab => wire_add_sub14_datab,
		result => wire_add_sub14_result
	  );
	wire_add_sub15_dataa <= ( slevel_w11c(55 DOWNTO 42));
	wire_add_sub15_datab <= ( wire_alt_sqrt_block2_w3560w & qlevel_w11c(1 DOWNTO 0));
	add_sub15 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		dataa => wire_add_sub15_dataa,
		datab => wire_add_sub15_datab,
		result => wire_add_sub15_result
	  );
	wire_add_sub16_dataa <= ( slevel_w12c(55 DOWNTO 41));
	wire_add_sub16_datab <= ( wire_rad_ff11c_w_lg_w_lg_w_lg_w_q_range3587w3590w3591w3592w & qlevel_w12c(1 DOWNTO 0));
	add_sub16 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 15
	  )
	  PORT MAP ( 
		dataa => wire_add_sub16_dataa,
		datab => wire_add_sub16_datab,
		result => wire_add_sub16_result
	  );
	wire_add_sub17_dataa <= ( slevel_w13c(55 DOWNTO 40));
	wire_add_sub17_datab <= ( wire_alt_sqrt_block2_w3622w & qlevel_w13c(1 DOWNTO 0));
	add_sub17 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 16
	  )
	  PORT MAP ( 
		dataa => wire_add_sub17_dataa,
		datab => wire_add_sub17_datab,
		result => wire_add_sub17_result
	  );
	wire_add_sub18_dataa <= ( slevel_w14c(55 DOWNTO 39));
	wire_add_sub18_datab <= ( wire_rad_ff13c_w_lg_w_lg_w_lg_w_q_range3649w3652w3653w3654w & qlevel_w14c(1 DOWNTO 0));
	add_sub18 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 17
	  )
	  PORT MAP ( 
		dataa => wire_add_sub18_dataa,
		datab => wire_add_sub18_datab,
		result => wire_add_sub18_result
	  );
	wire_add_sub19_dataa <= ( slevel_w15c(55 DOWNTO 38));
	wire_add_sub19_datab <= ( wire_alt_sqrt_block2_w3684w & qlevel_w15c(1 DOWNTO 0));
	add_sub19 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 18
	  )
	  PORT MAP ( 
		dataa => wire_add_sub19_dataa,
		datab => wire_add_sub19_datab,
		result => wire_add_sub19_result
	  );
	wire_add_sub20_dataa <= ( slevel_w16c(55 DOWNTO 37));
	wire_add_sub20_datab <= ( wire_rad_ff15c_w_lg_w_lg_w_lg_w_q_range3711w3714w3715w3716w & qlevel_w16c(1 DOWNTO 0));
	add_sub20 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 19
	  )
	  PORT MAP ( 
		dataa => wire_add_sub20_dataa,
		datab => wire_add_sub20_datab,
		result => wire_add_sub20_result
	  );
	wire_add_sub21_dataa <= ( slevel_w17c(55 DOWNTO 36));
	wire_add_sub21_datab <= ( wire_alt_sqrt_block2_w3746w & qlevel_w17c(1 DOWNTO 0));
	add_sub21 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 20
	  )
	  PORT MAP ( 
		dataa => wire_add_sub21_dataa,
		datab => wire_add_sub21_datab,
		result => wire_add_sub21_result
	  );
	wire_add_sub22_dataa <= ( slevel_w18c(55 DOWNTO 35));
	wire_add_sub22_datab <= ( wire_rad_ff17c_w_lg_w_lg_w_lg_w_q_range3773w3776w3777w3778w & qlevel_w18c(1 DOWNTO 0));
	add_sub22 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 21
	  )
	  PORT MAP ( 
		dataa => wire_add_sub22_dataa,
		datab => wire_add_sub22_datab,
		result => wire_add_sub22_result
	  );
	wire_add_sub23_dataa <= ( slevel_w19c(55 DOWNTO 34));
	wire_add_sub23_datab <= ( wire_alt_sqrt_block2_w3808w & qlevel_w19c(1 DOWNTO 0));
	add_sub23 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 22
	  )
	  PORT MAP ( 
		dataa => wire_add_sub23_dataa,
		datab => wire_add_sub23_datab,
		result => wire_add_sub23_result
	  );
	wire_add_sub24_dataa <= ( slevel_w20c(55 DOWNTO 33));
	wire_add_sub24_datab <= ( wire_rad_ff19c_w_lg_w_lg_w_lg_w_q_range3835w3838w3839w3840w & qlevel_w20c(1 DOWNTO 0));
	add_sub24 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 23
	  )
	  PORT MAP ( 
		dataa => wire_add_sub24_dataa,
		datab => wire_add_sub24_datab,
		result => wire_add_sub24_result
	  );
	wire_add_sub25_dataa <= ( slevel_w21c(55 DOWNTO 32));
	wire_add_sub25_datab <= ( wire_alt_sqrt_block2_w3870w & qlevel_w21c(1 DOWNTO 0));
	add_sub25 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 24
	  )
	  PORT MAP ( 
		dataa => wire_add_sub25_dataa,
		datab => wire_add_sub25_datab,
		result => wire_add_sub25_result
	  );
	wire_add_sub26_dataa <= ( slevel_w22c(55 DOWNTO 31));
	wire_add_sub26_datab <= ( wire_rad_ff21c_w_lg_w_lg_w_lg_w_q_range3897w3900w3901w3902w & qlevel_w22c(1 DOWNTO 0));
	add_sub26 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 25
	  )
	  PORT MAP ( 
		dataa => wire_add_sub26_dataa,
		datab => wire_add_sub26_datab,
		result => wire_add_sub26_result
	  );
	wire_add_sub27_dataa <= ( slevel_w23c(55 DOWNTO 30));
	wire_add_sub27_datab <= ( wire_alt_sqrt_block2_w3932w & qlevel_w23c(1 DOWNTO 0));
	add_sub27 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 26
	  )
	  PORT MAP ( 
		dataa => wire_add_sub27_dataa,
		datab => wire_add_sub27_datab,
		result => wire_add_sub27_result
	  );
	wire_add_sub28_dataa <= ( slevel_w24c(55 DOWNTO 29));
	wire_add_sub28_datab <= ( wire_rad_ff23c_w_lg_w_lg_w_lg_w_q_range3959w3962w3963w3964w & qlevel_w24c(1 DOWNTO 0));
	add_sub28 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 27
	  )
	  PORT MAP ( 
		dataa => wire_add_sub28_dataa,
		datab => wire_add_sub28_datab,
		result => wire_add_sub28_result
	  );
	wire_add_sub29_dataa <= ( slevel_w25c(55 DOWNTO 28));
	wire_add_sub29_datab <= ( wire_alt_sqrt_block2_w3994w & qlevel_w25c(1 DOWNTO 0));
	add_sub29 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 28
	  )
	  PORT MAP ( 
		dataa => wire_add_sub29_dataa,
		datab => wire_add_sub29_datab,
		result => wire_add_sub29_result
	  );
	wire_add_sub30_dataa <= ( slevel_w26c(55 DOWNTO 27));
	wire_add_sub30_datab <= ( wire_rad_ff25c_w_lg_w_lg_w_lg_w_q_range4020w4023w4024w4025w & qlevel_w26c(1 DOWNTO 0));
	add_sub30 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 29
	  )
	  PORT MAP ( 
		dataa => wire_add_sub30_dataa,
		datab => wire_add_sub30_datab,
		result => wire_add_sub30_result
	  );
	wire_add_sub31_dataa <= ( slevel_w27c(55 DOWNTO 28));
	wire_add_sub31_datab <= ( wire_alt_sqrt_block2_w4053w);
	add_sub31 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 28
	  )
	  PORT MAP ( 
		dataa => wire_add_sub31_dataa,
		datab => wire_add_sub31_datab,
		result => wire_add_sub31_result
	  );
	wire_add_sub32_dataa <= ( slevel_w28c(55 DOWNTO 28));
	wire_add_sub32_datab <= ( wire_rad_ff27c_w_lg_w_lg_w_lg_w_q_range4083w4086w4087w4088w);
	add_sub32 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 28
	  )
	  PORT MAP ( 
		dataa => wire_add_sub32_dataa,
		datab => wire_add_sub32_datab,
		result => wire_add_sub32_result
	  );
	wire_add_sub33_dataa <= ( slevel_w29c(55 DOWNTO 27));
	wire_add_sub33_datab <= ( wire_alt_sqrt_block2_w4126w);
	add_sub33 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 29
	  )
	  PORT MAP ( 
		dataa => wire_add_sub33_dataa,
		datab => wire_add_sub33_datab,
		result => wire_add_sub33_result
	  );
	wire_add_sub34_dataa <= ( slevel_w30c(55 DOWNTO 26));
	wire_add_sub34_datab <= ( wire_rad_ff29c_w_lg_w_lg_w_lg_w_q_range4160w4163w4164w4165w);
	add_sub34 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 30
	  )
	  PORT MAP ( 
		dataa => wire_add_sub34_dataa,
		datab => wire_add_sub34_datab,
		result => wire_add_sub34_result
	  );
	wire_add_sub35_dataa <= ( slevel_w31c(55 DOWNTO 25));
	wire_add_sub35_datab <= ( wire_alt_sqrt_block2_w4203w);
	add_sub35 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 31
	  )
	  PORT MAP ( 
		dataa => wire_add_sub35_dataa,
		datab => wire_add_sub35_datab,
		result => wire_add_sub35_result
	  );
	wire_add_sub36_dataa <= ( slevel_w32c(55 DOWNTO 24));
	wire_add_sub36_datab <= ( wire_rad_ff31c_w_lg_w_lg_w_lg_w_q_range4237w4240w4241w4242w);
	add_sub36 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 32
	  )
	  PORT MAP ( 
		dataa => wire_add_sub36_dataa,
		datab => wire_add_sub36_datab,
		result => wire_add_sub36_result
	  );
	wire_add_sub37_dataa <= ( slevel_w33c(55 DOWNTO 23));
	wire_add_sub37_datab <= ( wire_alt_sqrt_block2_w4280w);
	add_sub37 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 33
	  )
	  PORT MAP ( 
		dataa => wire_add_sub37_dataa,
		datab => wire_add_sub37_datab,
		result => wire_add_sub37_result
	  );
	wire_add_sub38_dataa <= ( slevel_w34c(55 DOWNTO 22));
	wire_add_sub38_datab <= ( wire_rad_ff33c_w_lg_w_lg_w_lg_w_q_range4314w4317w4318w4319w);
	add_sub38 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 34
	  )
	  PORT MAP ( 
		dataa => wire_add_sub38_dataa,
		datab => wire_add_sub38_datab,
		result => wire_add_sub38_result
	  );
	wire_add_sub39_dataa <= ( slevel_w35c(55 DOWNTO 21));
	wire_add_sub39_datab <= ( wire_alt_sqrt_block2_w4357w);
	add_sub39 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 35
	  )
	  PORT MAP ( 
		dataa => wire_add_sub39_dataa,
		datab => wire_add_sub39_datab,
		result => wire_add_sub39_result
	  );
	wire_add_sub4_dataa <= ( slevel_w0c(55 DOWNTO 53));
	wire_add_sub4_datab <= ( qlevel_w0c(2 DOWNTO 0));
	add_sub4 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 3
	  )
	  PORT MAP ( 
		dataa => wire_add_sub4_dataa,
		datab => wire_add_sub4_datab,
		result => wire_add_sub4_result
	  );
	wire_add_sub40_dataa <= ( slevel_w36c(55 DOWNTO 20));
	wire_add_sub40_datab <= ( wire_rad_ff35c_w_lg_w_lg_w_lg_w_q_range4391w4394w4395w4396w);
	add_sub40 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 36
	  )
	  PORT MAP ( 
		dataa => wire_add_sub40_dataa,
		datab => wire_add_sub40_datab,
		result => wire_add_sub40_result
	  );
	wire_add_sub41_dataa <= ( slevel_w37c(55 DOWNTO 19));
	wire_add_sub41_datab <= ( wire_alt_sqrt_block2_w4434w);
	add_sub41 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 37
	  )
	  PORT MAP ( 
		dataa => wire_add_sub41_dataa,
		datab => wire_add_sub41_datab,
		result => wire_add_sub41_result
	  );
	wire_add_sub42_dataa <= ( slevel_w38c(55 DOWNTO 18));
	wire_add_sub42_datab <= ( wire_rad_ff37c_w_lg_w_lg_w_lg_w_q_range4468w4471w4472w4473w);
	add_sub42 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 38
	  )
	  PORT MAP ( 
		dataa => wire_add_sub42_dataa,
		datab => wire_add_sub42_datab,
		result => wire_add_sub42_result
	  );
	wire_add_sub43_dataa <= ( slevel_w39c(55 DOWNTO 17));
	wire_add_sub43_datab <= ( wire_alt_sqrt_block2_w4511w);
	add_sub43 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 39
	  )
	  PORT MAP ( 
		dataa => wire_add_sub43_dataa,
		datab => wire_add_sub43_datab,
		result => wire_add_sub43_result
	  );
	wire_add_sub44_dataa <= ( slevel_w40c(55 DOWNTO 16));
	wire_add_sub44_datab <= ( wire_rad_ff39c_w_lg_w_lg_w_lg_w_q_range4545w4548w4549w4550w);
	add_sub44 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 40
	  )
	  PORT MAP ( 
		dataa => wire_add_sub44_dataa,
		datab => wire_add_sub44_datab,
		result => wire_add_sub44_result
	  );
	wire_add_sub45_dataa <= ( slevel_w41c(55 DOWNTO 15));
	wire_add_sub45_datab <= ( wire_alt_sqrt_block2_w4588w);
	add_sub45 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 41
	  )
	  PORT MAP ( 
		dataa => wire_add_sub45_dataa,
		datab => wire_add_sub45_datab,
		result => wire_add_sub45_result
	  );
	wire_add_sub46_dataa <= ( slevel_w42c(55 DOWNTO 14));
	wire_add_sub46_datab <= ( wire_rad_ff41c_w_lg_w_lg_w_lg_w_q_range4622w4625w4626w4627w);
	add_sub46 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 42
	  )
	  PORT MAP ( 
		dataa => wire_add_sub46_dataa,
		datab => wire_add_sub46_datab,
		result => wire_add_sub46_result
	  );
	wire_add_sub47_dataa <= ( slevel_w43c(55 DOWNTO 13));
	wire_add_sub47_datab <= ( wire_alt_sqrt_block2_w4665w);
	add_sub47 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 43
	  )
	  PORT MAP ( 
		dataa => wire_add_sub47_dataa,
		datab => wire_add_sub47_datab,
		result => wire_add_sub47_result
	  );
	wire_add_sub48_dataa <= ( slevel_w44c(55 DOWNTO 12));
	wire_add_sub48_datab <= ( wire_rad_ff43c_w_lg_w_lg_w_lg_w_q_range4699w4702w4703w4704w);
	add_sub48 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 44
	  )
	  PORT MAP ( 
		dataa => wire_add_sub48_dataa,
		datab => wire_add_sub48_datab,
		result => wire_add_sub48_result
	  );
	wire_add_sub49_dataa <= ( slevel_w45c(55 DOWNTO 11));
	wire_add_sub49_datab <= ( wire_alt_sqrt_block2_w4742w);
	add_sub49 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 45
	  )
	  PORT MAP ( 
		dataa => wire_add_sub49_dataa,
		datab => wire_add_sub49_datab,
		result => wire_add_sub49_result
	  );
	wire_add_sub5_dataa <= ( slevel_w1c(55 DOWNTO 52));
	wire_add_sub5_datab <= ( qlevel_w1c(3 DOWNTO 0));
	add_sub5 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 4
	  )
	  PORT MAP ( 
		dataa => wire_add_sub5_dataa,
		datab => wire_add_sub5_datab,
		result => wire_add_sub5_result
	  );
	wire_add_sub50_dataa <= ( slevel_w46c(55 DOWNTO 10));
	wire_add_sub50_datab <= ( wire_rad_ff45c_w_lg_w_lg_w_lg_w_q_range4776w4779w4780w4781w);
	add_sub50 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 46
	  )
	  PORT MAP ( 
		dataa => wire_add_sub50_dataa,
		datab => wire_add_sub50_datab,
		result => wire_add_sub50_result
	  );
	wire_add_sub51_dataa <= ( slevel_w47c(55 DOWNTO 9));
	wire_add_sub51_datab <= ( wire_alt_sqrt_block2_w4819w);
	add_sub51 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 47
	  )
	  PORT MAP ( 
		dataa => wire_add_sub51_dataa,
		datab => wire_add_sub51_datab,
		result => wire_add_sub51_result
	  );
	wire_add_sub52_dataa <= ( slevel_w48c(55 DOWNTO 8));
	wire_add_sub52_datab <= ( wire_rad_ff47c_w_lg_w_lg_w_lg_w_q_range4853w4856w4857w4858w);
	add_sub52 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 48
	  )
	  PORT MAP ( 
		dataa => wire_add_sub52_dataa,
		datab => wire_add_sub52_datab,
		result => wire_add_sub52_result
	  );
	wire_add_sub53_dataa <= ( slevel_w49c(55 DOWNTO 7));
	wire_add_sub53_datab <= ( wire_alt_sqrt_block2_w4896w);
	add_sub53 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 49
	  )
	  PORT MAP ( 
		dataa => wire_add_sub53_dataa,
		datab => wire_add_sub53_datab,
		result => wire_add_sub53_result
	  );
	wire_add_sub54_dataa <= ( slevel_w50c(55 DOWNTO 6));
	wire_add_sub54_datab <= ( wire_rad_ff49c_w_lg_w_lg_w_lg_w_q_range4930w4933w4934w4935w);
	add_sub54 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 50
	  )
	  PORT MAP ( 
		dataa => wire_add_sub54_dataa,
		datab => wire_add_sub54_datab,
		result => wire_add_sub54_result
	  );
	wire_add_sub55_dataa <= ( slevel_w51c(55 DOWNTO 5));
	wire_add_sub55_datab <= ( wire_alt_sqrt_block2_w4973w);
	add_sub55 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 51
	  )
	  PORT MAP ( 
		dataa => wire_add_sub55_dataa,
		datab => wire_add_sub55_datab,
		result => wire_add_sub55_result
	  );
	wire_add_sub56_dataa <= ( slevel_w52c(55 DOWNTO 4));
	wire_add_sub56_datab <= ( wire_rad_ff51c_w_lg_w_lg_w_lg_w_q_range5007w5010w5011w5012w);
	add_sub56 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 52
	  )
	  PORT MAP ( 
		dataa => wire_add_sub56_dataa,
		datab => wire_add_sub56_datab,
		result => wire_add_sub56_result
	  );
	wire_add_sub57_dataa <= ( slevel_w53c(55 DOWNTO 3));
	wire_add_sub57_datab <= ( qlevel_w53c(55 DOWNTO 54) & wire_alt_sqrt_block2_w5051w);
	add_sub57 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 53
	  )
	  PORT MAP ( 
		dataa => wire_add_sub57_dataa,
		datab => wire_add_sub57_datab,
		result => wire_add_sub57_result
	  );
	wire_add_sub6_dataa <= ( slevel_w2c(55 DOWNTO 51));
	wire_add_sub6_datab <= ( wire_rad_ff1c_w_lg_w_lg_w_lg_w_q_range3277w3280w3281w3282w & qlevel_w2c(1 DOWNTO 0));
	add_sub6 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 5
	  )
	  PORT MAP ( 
		dataa => wire_add_sub6_dataa,
		datab => wire_add_sub6_datab,
		result => wire_add_sub6_result
	  );
	wire_add_sub7_dataa <= ( slevel_w3c(55 DOWNTO 50));
	wire_add_sub7_datab <= ( wire_alt_sqrt_block2_w3312w & qlevel_w3c(1 DOWNTO 0));
	add_sub7 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 6
	  )
	  PORT MAP ( 
		dataa => wire_add_sub7_dataa,
		datab => wire_add_sub7_datab,
		result => wire_add_sub7_result
	  );
	wire_add_sub8_dataa <= ( slevel_w4c(55 DOWNTO 49));
	wire_add_sub8_datab <= ( wire_rad_ff3c_w_lg_w_lg_w_lg_w_q_range3339w3342w3343w3344w & qlevel_w4c(1 DOWNTO 0));
	add_sub8 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 7
	  )
	  PORT MAP ( 
		dataa => wire_add_sub8_dataa,
		datab => wire_add_sub8_datab,
		result => wire_add_sub8_result
	  );
	wire_add_sub9_dataa <= ( slevel_w5c(55 DOWNTO 48));
	wire_add_sub9_datab <= ( wire_alt_sqrt_block2_w3374w & qlevel_w5c(1 DOWNTO 0));
	add_sub9 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 8
	  )
	  PORT MAP ( 
		dataa => wire_add_sub9_dataa,
		datab => wire_add_sub9_datab,
		result => wire_add_sub9_result
	  );

 END RTL; --fp_sqrt_dp_alt_sqrt_block_kgb

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 56 reg 2983 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  fp_sqrt_dp_altfp_sqrt_lqd IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clk_en	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC;
		 data	:	IN  STD_LOGIC_VECTOR (63 DOWNTO 0);
		 result	:	OUT  STD_LOGIC_VECTOR (63 DOWNTO 0)
	 ); 
 END fp_sqrt_dp_altfp_sqrt_lqd;

 ARCHITECTURE RTL OF fp_sqrt_dp_altfp_sqrt_lqd IS

	 SIGNAL  wire_alt_sqrt_block2_root_result	:	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL	 exp_all_one_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff1	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff20c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff210c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff211c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff212c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff213c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff214c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff215c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff216c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff217c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff218c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff219c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff21c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff220c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff221c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff222c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff223c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff224c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff225c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff226c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff22c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff23c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff24c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff25c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff26c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff27c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff28c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_ff29c	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_in_ff	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range78w82w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range33w37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range38w42w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range43w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range48w52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range53w57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range58w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range63w67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range68w72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range73w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range78w80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range33w35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range38w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range43w45w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range48w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range53w55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range58w60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range63w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range68w70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_lg_w_q_range73w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range43w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range68w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_exp_in_ff_w_q_range73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exp_not_zero_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_result_ff	:	STD_LOGIC_VECTOR(10 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff25	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 infinity_ff26	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_in_ff	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range83w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range269w270w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range271w272w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range236w276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_lg_w_q_range271w272w273w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range113w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range116w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range119w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range122w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range125w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range128w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range131w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range134w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range137w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range140w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range86w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range143w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range146w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range149w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range152w154w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range155w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range158w160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range161w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range164w166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range167w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range170w172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range89w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range173w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range176w178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range179w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range182w184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range185w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range188w190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range191w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range194w196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range197w199w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range200w202w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range92w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range203w205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range206w208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range209w211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range212w214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range215w217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range218w220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range221w223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range224w226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range227w229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range230w232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range95w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range233w235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range236w238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range98w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range101w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range104w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range107w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_lg_w_q_range110w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range83w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range86w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range152w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range200w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range269w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range271w	:	STD_LOGIC_VECTOR (50 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_man_in_ff_w_q_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_not_zero_ff	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_not_zero_ff_w_lg_q239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_result_ff	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_rounding_ff	:	STD_LOGIC_VECTOR(51 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_rounding_ff_w_lg_q285w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_man_rounding_ff_w_lg_w_lg_q285w286w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL	 nan_man_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff25	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 nan_man_ff26	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_sign_node_ff_w_lg_q244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 sign_node_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff25	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff26	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff27	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff28	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_node_ff29	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff0	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff1	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff2	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff3	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff4	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff5	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff6	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff7	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff8	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff9	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff10	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff11	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff12	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff13	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff14	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff15	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff16	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff17	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff18	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff19	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff20	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff21	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff22	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff23	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff24	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff25	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 zero_exp_ff26	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub1_dataa	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub1_datab	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub1_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_add_sub3_datab	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_add_sub3_result	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_ff2_w260w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_preadjust_w268w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_ff2_w260w261w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_exp_ff2_w260w261w262w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_lg_preadjust_w277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  bias :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_all_one_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_div_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_ff2_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  exp_not_zero_w :	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  infinitycondition_w :	STD_LOGIC;
	 SIGNAL  man_not_zero_w :	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  man_root_result_w :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  nancondition_w :	STD_LOGIC;
	 SIGNAL  preadjust_w :	STD_LOGIC;
	 SIGNAL  radicand_w :	STD_LOGIC_VECTOR (54 DOWNTO 0);
	 SIGNAL  roundbit_w :	STD_LOGIC;
	 SIGNAL  wire_w_data_range27w	:	STD_LOGIC_VECTOR (51 DOWNTO 0);
	 SIGNAL  wire_w_data_range26w	:	STD_LOGIC_VECTOR (10 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range41w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range66w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_all_one_w_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_not_zero_w_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range84w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range198w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_not_zero_w_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  fp_sqrt_dp_alt_sqrt_block_kgb
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		rad	:	IN  STD_LOGIC_VECTOR(54 DOWNTO 0);
		root_result	:	OUT  STD_LOGIC_VECTOR(53 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	loop208 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_exp_ff2_w260w(i) <= exp_ff2_w(i) AND zero_exp_ff26;
	END GENERATE loop208;
	wire_w_lg_preadjust_w268w(0) <= NOT preadjust_w;
	loop209 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_exp_ff2_w260w261w(i) <= wire_w_lg_exp_ff2_w260w(i) OR nan_man_ff26;
	END GENERATE loop209;
	loop210 : FOR i IN 0 TO 10 GENERATE 
		wire_w_lg_w_lg_w_lg_exp_ff2_w260w261w262w(i) <= wire_w_lg_w_lg_exp_ff2_w260w261w(i) OR infinity_ff26;
	END GENERATE loop210;
	wire_w_lg_preadjust_w277w(0) <= preadjust_w OR wire_man_in_ff_w_lg_w_q_range236w276w(0);
	bias <= ( "0" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1" & "1");
	exp_all_one_w <= ( wire_exp_in_ff_w_lg_w_q_range78w82w & wire_exp_in_ff_w_lg_w_q_range73w77w & wire_exp_in_ff_w_lg_w_q_range68w72w & wire_exp_in_ff_w_lg_w_q_range63w67w & wire_exp_in_ff_w_lg_w_q_range58w62w & wire_exp_in_ff_w_lg_w_q_range53w57w & wire_exp_in_ff_w_lg_w_q_range48w52w & wire_exp_in_ff_w_lg_w_q_range43w47w & wire_exp_in_ff_w_lg_w_q_range38w42w & wire_exp_in_ff_w_lg_w_q_range33w37w & exp_in_ff(0));
	exp_div_w <= ( wire_add_sub1_result(11 DOWNTO 1));
	exp_ff2_w <= exp_ff226c;
	exp_not_zero_w <= ( wire_exp_in_ff_w_lg_w_q_range78w80w & wire_exp_in_ff_w_lg_w_q_range73w75w & wire_exp_in_ff_w_lg_w_q_range68w70w & wire_exp_in_ff_w_lg_w_q_range63w65w & wire_exp_in_ff_w_lg_w_q_range58w60w & wire_exp_in_ff_w_lg_w_q_range53w55w & wire_exp_in_ff_w_lg_w_q_range48w50w & wire_exp_in_ff_w_lg_w_q_range43w45w & wire_exp_in_ff_w_lg_w_q_range38w40w & wire_exp_in_ff_w_lg_w_q_range33w35w & exp_in_ff(0));
	infinitycondition_w <= (wire_man_not_zero_ff_w_lg_q239w(0) AND exp_all_one_ff);
	man_not_zero_w <= ( wire_man_in_ff_w_lg_w_q_range236w238w & wire_man_in_ff_w_lg_w_q_range233w235w & wire_man_in_ff_w_lg_w_q_range230w232w & wire_man_in_ff_w_lg_w_q_range227w229w & wire_man_in_ff_w_lg_w_q_range224w226w & wire_man_in_ff_w_lg_w_q_range221w223w & wire_man_in_ff_w_lg_w_q_range218w220w & wire_man_in_ff_w_lg_w_q_range215w217w & wire_man_in_ff_w_lg_w_q_range212w214w & wire_man_in_ff_w_lg_w_q_range209w211w & wire_man_in_ff_w_lg_w_q_range206w208w & wire_man_in_ff_w_lg_w_q_range203w205w & wire_man_in_ff_w_lg_w_q_range200w202w & wire_man_in_ff_w_lg_w_q_range197w199w & wire_man_in_ff_w_lg_w_q_range194w196w & wire_man_in_ff_w_lg_w_q_range191w193w & wire_man_in_ff_w_lg_w_q_range188w190w & wire_man_in_ff_w_lg_w_q_range185w187w & wire_man_in_ff_w_lg_w_q_range182w184w & wire_man_in_ff_w_lg_w_q_range179w181w & wire_man_in_ff_w_lg_w_q_range176w178w & wire_man_in_ff_w_lg_w_q_range173w175w & wire_man_in_ff_w_lg_w_q_range170w172w & wire_man_in_ff_w_lg_w_q_range167w169w & wire_man_in_ff_w_lg_w_q_range164w166w & wire_man_in_ff_w_lg_w_q_range161w163w & wire_man_in_ff_w_lg_w_q_range158w160w & wire_man_in_ff_w_lg_w_q_range155w157w & wire_man_in_ff_w_lg_w_q_range152w154w & wire_man_in_ff_w_lg_w_q_range149w151w & wire_man_in_ff_w_lg_w_q_range146w148w & wire_man_in_ff_w_lg_w_q_range143w145w & wire_man_in_ff_w_lg_w_q_range140w142w & wire_man_in_ff_w_lg_w_q_range137w139w & wire_man_in_ff_w_lg_w_q_range134w136w & wire_man_in_ff_w_lg_w_q_range131w133w & wire_man_in_ff_w_lg_w_q_range128w130w & wire_man_in_ff_w_lg_w_q_range125w127w & wire_man_in_ff_w_lg_w_q_range122w124w & wire_man_in_ff_w_lg_w_q_range119w121w & wire_man_in_ff_w_lg_w_q_range116w118w & wire_man_in_ff_w_lg_w_q_range113w115w & wire_man_in_ff_w_lg_w_q_range110w112w & wire_man_in_ff_w_lg_w_q_range107w109w & wire_man_in_ff_w_lg_w_q_range104w106w & wire_man_in_ff_w_lg_w_q_range101w103w & wire_man_in_ff_w_lg_w_q_range98w100w & wire_man_in_ff_w_lg_w_q_range95w97w & wire_man_in_ff_w_lg_w_q_range92w94w & wire_man_in_ff_w_lg_w_q_range89w91w & wire_man_in_ff_w_lg_w_q_range86w88w
 & man_in_ff(0));
	man_root_result_w <= wire_alt_sqrt_block2_root_result;
	nancondition_w <= ((sign_node_ff1 AND exp_not_zero_ff) OR (exp_all_one_ff AND man_not_zero_ff));
	preadjust_w <= exp_in_ff(0);
	radicand_w <= ( wire_w_lg_preadjust_w268w & wire_w_lg_preadjust_w277w & wire_man_in_ff_w_lg_w_lg_w_q_range271w272w273w & wire_man_in_ff_w_lg_w_q_range83w267w & "0");
	result <= ( sign_node_ff29 & exp_result_ff & man_result_ff);
	roundbit_w <= wire_alt_sqrt_block2_root_result(0);
	wire_w_data_range27w <= data(51 DOWNTO 0);
	wire_w_data_range26w <= data(62 DOWNTO 52);
	wire_w_exp_all_one_w_range31w(0) <= exp_all_one_w(0);
	wire_w_exp_all_one_w_range36w(0) <= exp_all_one_w(1);
	wire_w_exp_all_one_w_range41w(0) <= exp_all_one_w(2);
	wire_w_exp_all_one_w_range46w(0) <= exp_all_one_w(3);
	wire_w_exp_all_one_w_range51w(0) <= exp_all_one_w(4);
	wire_w_exp_all_one_w_range56w(0) <= exp_all_one_w(5);
	wire_w_exp_all_one_w_range61w(0) <= exp_all_one_w(6);
	wire_w_exp_all_one_w_range66w(0) <= exp_all_one_w(7);
	wire_w_exp_all_one_w_range71w(0) <= exp_all_one_w(8);
	wire_w_exp_all_one_w_range76w(0) <= exp_all_one_w(9);
	wire_w_exp_not_zero_w_range29w(0) <= exp_not_zero_w(0);
	wire_w_exp_not_zero_w_range34w(0) <= exp_not_zero_w(1);
	wire_w_exp_not_zero_w_range39w(0) <= exp_not_zero_w(2);
	wire_w_exp_not_zero_w_range44w(0) <= exp_not_zero_w(3);
	wire_w_exp_not_zero_w_range49w(0) <= exp_not_zero_w(4);
	wire_w_exp_not_zero_w_range54w(0) <= exp_not_zero_w(5);
	wire_w_exp_not_zero_w_range59w(0) <= exp_not_zero_w(6);
	wire_w_exp_not_zero_w_range64w(0) <= exp_not_zero_w(7);
	wire_w_exp_not_zero_w_range69w(0) <= exp_not_zero_w(8);
	wire_w_exp_not_zero_w_range74w(0) <= exp_not_zero_w(9);
	wire_w_man_not_zero_w_range84w(0) <= man_not_zero_w(0);
	wire_w_man_not_zero_w_range114w(0) <= man_not_zero_w(10);
	wire_w_man_not_zero_w_range117w(0) <= man_not_zero_w(11);
	wire_w_man_not_zero_w_range120w(0) <= man_not_zero_w(12);
	wire_w_man_not_zero_w_range123w(0) <= man_not_zero_w(13);
	wire_w_man_not_zero_w_range126w(0) <= man_not_zero_w(14);
	wire_w_man_not_zero_w_range129w(0) <= man_not_zero_w(15);
	wire_w_man_not_zero_w_range132w(0) <= man_not_zero_w(16);
	wire_w_man_not_zero_w_range135w(0) <= man_not_zero_w(17);
	wire_w_man_not_zero_w_range138w(0) <= man_not_zero_w(18);
	wire_w_man_not_zero_w_range141w(0) <= man_not_zero_w(19);
	wire_w_man_not_zero_w_range87w(0) <= man_not_zero_w(1);
	wire_w_man_not_zero_w_range144w(0) <= man_not_zero_w(20);
	wire_w_man_not_zero_w_range147w(0) <= man_not_zero_w(21);
	wire_w_man_not_zero_w_range150w(0) <= man_not_zero_w(22);
	wire_w_man_not_zero_w_range153w(0) <= man_not_zero_w(23);
	wire_w_man_not_zero_w_range156w(0) <= man_not_zero_w(24);
	wire_w_man_not_zero_w_range159w(0) <= man_not_zero_w(25);
	wire_w_man_not_zero_w_range162w(0) <= man_not_zero_w(26);
	wire_w_man_not_zero_w_range165w(0) <= man_not_zero_w(27);
	wire_w_man_not_zero_w_range168w(0) <= man_not_zero_w(28);
	wire_w_man_not_zero_w_range171w(0) <= man_not_zero_w(29);
	wire_w_man_not_zero_w_range90w(0) <= man_not_zero_w(2);
	wire_w_man_not_zero_w_range174w(0) <= man_not_zero_w(30);
	wire_w_man_not_zero_w_range177w(0) <= man_not_zero_w(31);
	wire_w_man_not_zero_w_range180w(0) <= man_not_zero_w(32);
	wire_w_man_not_zero_w_range183w(0) <= man_not_zero_w(33);
	wire_w_man_not_zero_w_range186w(0) <= man_not_zero_w(34);
	wire_w_man_not_zero_w_range189w(0) <= man_not_zero_w(35);
	wire_w_man_not_zero_w_range192w(0) <= man_not_zero_w(36);
	wire_w_man_not_zero_w_range195w(0) <= man_not_zero_w(37);
	wire_w_man_not_zero_w_range198w(0) <= man_not_zero_w(38);
	wire_w_man_not_zero_w_range201w(0) <= man_not_zero_w(39);
	wire_w_man_not_zero_w_range93w(0) <= man_not_zero_w(3);
	wire_w_man_not_zero_w_range204w(0) <= man_not_zero_w(40);
	wire_w_man_not_zero_w_range207w(0) <= man_not_zero_w(41);
	wire_w_man_not_zero_w_range210w(0) <= man_not_zero_w(42);
	wire_w_man_not_zero_w_range213w(0) <= man_not_zero_w(43);
	wire_w_man_not_zero_w_range216w(0) <= man_not_zero_w(44);
	wire_w_man_not_zero_w_range219w(0) <= man_not_zero_w(45);
	wire_w_man_not_zero_w_range222w(0) <= man_not_zero_w(46);
	wire_w_man_not_zero_w_range225w(0) <= man_not_zero_w(47);
	wire_w_man_not_zero_w_range228w(0) <= man_not_zero_w(48);
	wire_w_man_not_zero_w_range231w(0) <= man_not_zero_w(49);
	wire_w_man_not_zero_w_range96w(0) <= man_not_zero_w(4);
	wire_w_man_not_zero_w_range234w(0) <= man_not_zero_w(50);
	wire_w_man_not_zero_w_range99w(0) <= man_not_zero_w(5);
	wire_w_man_not_zero_w_range102w(0) <= man_not_zero_w(6);
	wire_w_man_not_zero_w_range105w(0) <= man_not_zero_w(7);
	wire_w_man_not_zero_w_range108w(0) <= man_not_zero_w(8);
	wire_w_man_not_zero_w_range111w(0) <= man_not_zero_w(9);
	alt_sqrt_block2 :  fp_sqrt_dp_alt_sqrt_block_kgb
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		rad => radicand_w,
		root_result => wire_alt_sqrt_block2_root_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_all_one_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_all_one_ff <= exp_all_one_w(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff1 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff1 <= exp_div_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff20c <= exp_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff210c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff210c <= exp_ff29c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff211c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff211c <= exp_ff210c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff212c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff212c <= exp_ff211c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff213c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff213c <= exp_ff212c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff214c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff214c <= exp_ff213c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff215c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff215c <= exp_ff214c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff216c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff216c <= exp_ff215c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff217c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff217c <= exp_ff216c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff218c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff218c <= exp_ff217c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff219c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff219c <= exp_ff218c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff21c <= exp_ff20c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff220c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff220c <= exp_ff219c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff221c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff221c <= exp_ff220c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff222c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff222c <= exp_ff221c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff223c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff223c <= exp_ff222c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff224c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff224c <= exp_ff223c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff225c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff225c <= exp_ff224c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff226c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff226c <= exp_ff225c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff22c <= exp_ff21c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff23c <= exp_ff22c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff24c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff24c <= exp_ff23c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff25c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff25c <= exp_ff24c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff26c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff26c <= exp_ff25c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff27c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff27c <= exp_ff26c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff28c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff28c <= exp_ff27c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_ff29c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_ff29c <= exp_ff28c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_in_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_in_ff <= wire_w_data_range26w;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_in_ff_w_lg_w_q_range78w82w(0) <= wire_exp_in_ff_w_q_range78w(0) AND wire_w_exp_all_one_w_range76w(0);
	wire_exp_in_ff_w_lg_w_q_range33w37w(0) <= wire_exp_in_ff_w_q_range33w(0) AND wire_w_exp_all_one_w_range31w(0);
	wire_exp_in_ff_w_lg_w_q_range38w42w(0) <= wire_exp_in_ff_w_q_range38w(0) AND wire_w_exp_all_one_w_range36w(0);
	wire_exp_in_ff_w_lg_w_q_range43w47w(0) <= wire_exp_in_ff_w_q_range43w(0) AND wire_w_exp_all_one_w_range41w(0);
	wire_exp_in_ff_w_lg_w_q_range48w52w(0) <= wire_exp_in_ff_w_q_range48w(0) AND wire_w_exp_all_one_w_range46w(0);
	wire_exp_in_ff_w_lg_w_q_range53w57w(0) <= wire_exp_in_ff_w_q_range53w(0) AND wire_w_exp_all_one_w_range51w(0);
	wire_exp_in_ff_w_lg_w_q_range58w62w(0) <= wire_exp_in_ff_w_q_range58w(0) AND wire_w_exp_all_one_w_range56w(0);
	wire_exp_in_ff_w_lg_w_q_range63w67w(0) <= wire_exp_in_ff_w_q_range63w(0) AND wire_w_exp_all_one_w_range61w(0);
	wire_exp_in_ff_w_lg_w_q_range68w72w(0) <= wire_exp_in_ff_w_q_range68w(0) AND wire_w_exp_all_one_w_range66w(0);
	wire_exp_in_ff_w_lg_w_q_range73w77w(0) <= wire_exp_in_ff_w_q_range73w(0) AND wire_w_exp_all_one_w_range71w(0);
	wire_exp_in_ff_w_lg_w_q_range78w80w(0) <= wire_exp_in_ff_w_q_range78w(0) OR wire_w_exp_not_zero_w_range74w(0);
	wire_exp_in_ff_w_lg_w_q_range33w35w(0) <= wire_exp_in_ff_w_q_range33w(0) OR wire_w_exp_not_zero_w_range29w(0);
	wire_exp_in_ff_w_lg_w_q_range38w40w(0) <= wire_exp_in_ff_w_q_range38w(0) OR wire_w_exp_not_zero_w_range34w(0);
	wire_exp_in_ff_w_lg_w_q_range43w45w(0) <= wire_exp_in_ff_w_q_range43w(0) OR wire_w_exp_not_zero_w_range39w(0);
	wire_exp_in_ff_w_lg_w_q_range48w50w(0) <= wire_exp_in_ff_w_q_range48w(0) OR wire_w_exp_not_zero_w_range44w(0);
	wire_exp_in_ff_w_lg_w_q_range53w55w(0) <= wire_exp_in_ff_w_q_range53w(0) OR wire_w_exp_not_zero_w_range49w(0);
	wire_exp_in_ff_w_lg_w_q_range58w60w(0) <= wire_exp_in_ff_w_q_range58w(0) OR wire_w_exp_not_zero_w_range54w(0);
	wire_exp_in_ff_w_lg_w_q_range63w65w(0) <= wire_exp_in_ff_w_q_range63w(0) OR wire_w_exp_not_zero_w_range59w(0);
	wire_exp_in_ff_w_lg_w_q_range68w70w(0) <= wire_exp_in_ff_w_q_range68w(0) OR wire_w_exp_not_zero_w_range64w(0);
	wire_exp_in_ff_w_lg_w_q_range73w75w(0) <= wire_exp_in_ff_w_q_range73w(0) OR wire_w_exp_not_zero_w_range69w(0);
	wire_exp_in_ff_w_q_range78w(0) <= exp_in_ff(10);
	wire_exp_in_ff_w_q_range33w(0) <= exp_in_ff(1);
	wire_exp_in_ff_w_q_range38w(0) <= exp_in_ff(2);
	wire_exp_in_ff_w_q_range43w(0) <= exp_in_ff(3);
	wire_exp_in_ff_w_q_range48w(0) <= exp_in_ff(4);
	wire_exp_in_ff_w_q_range53w(0) <= exp_in_ff(5);
	wire_exp_in_ff_w_q_range58w(0) <= exp_in_ff(6);
	wire_exp_in_ff_w_q_range63w(0) <= exp_in_ff(7);
	wire_exp_in_ff_w_q_range68w(0) <= exp_in_ff(8);
	wire_exp_in_ff_w_q_range73w(0) <= exp_in_ff(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_not_zero_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_not_zero_ff <= exp_not_zero_w(10);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_result_ff <= wire_w_lg_w_lg_w_lg_exp_ff2_w260w261w262w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff0 <= (infinitycondition_w AND wire_sign_node_ff_w_lg_q244w(0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff1 <= infinity_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff2 <= infinity_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff3 <= infinity_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff4 <= infinity_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff5 <= infinity_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff6 <= infinity_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff7 <= infinity_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff8 <= infinity_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff9 <= infinity_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff10 <= infinity_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff11 <= infinity_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff12 <= infinity_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff13 <= infinity_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff14 <= infinity_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff15 <= infinity_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff16 <= infinity_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff17 <= infinity_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff18 <= infinity_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff19 <= infinity_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff20 <= infinity_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff21 <= infinity_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff22 <= infinity_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff23 <= infinity_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff24 <= infinity_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff25 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff25 <= infinity_ff24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN infinity_ff26 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN infinity_ff26 <= infinity_ff25;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_in_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_in_ff <= wire_w_data_range27w;
			END IF;
		END IF;
	END PROCESS;
	wire_man_in_ff_w_lg_w_q_range83w267w(0) <= wire_man_in_ff_w_q_range83w(0) AND preadjust_w;
	loop211 : FOR i IN 0 TO 50 GENERATE 
		wire_man_in_ff_w_lg_w_q_range269w270w(i) <= wire_man_in_ff_w_q_range269w(i) AND wire_w_lg_preadjust_w268w(0);
	END GENERATE loop211;
	loop212 : FOR i IN 0 TO 50 GENERATE 
		wire_man_in_ff_w_lg_w_q_range271w272w(i) <= wire_man_in_ff_w_q_range271w(i) AND preadjust_w;
	END GENERATE loop212;
	wire_man_in_ff_w_lg_w_q_range236w276w(0) <= wire_man_in_ff_w_q_range236w(0) AND wire_w_lg_preadjust_w268w(0);
	loop213 : FOR i IN 0 TO 50 GENERATE 
		wire_man_in_ff_w_lg_w_lg_w_q_range271w272w273w(i) <= wire_man_in_ff_w_lg_w_q_range271w272w(i) OR wire_man_in_ff_w_lg_w_q_range269w270w(i);
	END GENERATE loop213;
	wire_man_in_ff_w_lg_w_q_range113w115w(0) <= wire_man_in_ff_w_q_range113w(0) OR wire_w_man_not_zero_w_range111w(0);
	wire_man_in_ff_w_lg_w_q_range116w118w(0) <= wire_man_in_ff_w_q_range116w(0) OR wire_w_man_not_zero_w_range114w(0);
	wire_man_in_ff_w_lg_w_q_range119w121w(0) <= wire_man_in_ff_w_q_range119w(0) OR wire_w_man_not_zero_w_range117w(0);
	wire_man_in_ff_w_lg_w_q_range122w124w(0) <= wire_man_in_ff_w_q_range122w(0) OR wire_w_man_not_zero_w_range120w(0);
	wire_man_in_ff_w_lg_w_q_range125w127w(0) <= wire_man_in_ff_w_q_range125w(0) OR wire_w_man_not_zero_w_range123w(0);
	wire_man_in_ff_w_lg_w_q_range128w130w(0) <= wire_man_in_ff_w_q_range128w(0) OR wire_w_man_not_zero_w_range126w(0);
	wire_man_in_ff_w_lg_w_q_range131w133w(0) <= wire_man_in_ff_w_q_range131w(0) OR wire_w_man_not_zero_w_range129w(0);
	wire_man_in_ff_w_lg_w_q_range134w136w(0) <= wire_man_in_ff_w_q_range134w(0) OR wire_w_man_not_zero_w_range132w(0);
	wire_man_in_ff_w_lg_w_q_range137w139w(0) <= wire_man_in_ff_w_q_range137w(0) OR wire_w_man_not_zero_w_range135w(0);
	wire_man_in_ff_w_lg_w_q_range140w142w(0) <= wire_man_in_ff_w_q_range140w(0) OR wire_w_man_not_zero_w_range138w(0);
	wire_man_in_ff_w_lg_w_q_range86w88w(0) <= wire_man_in_ff_w_q_range86w(0) OR wire_w_man_not_zero_w_range84w(0);
	wire_man_in_ff_w_lg_w_q_range143w145w(0) <= wire_man_in_ff_w_q_range143w(0) OR wire_w_man_not_zero_w_range141w(0);
	wire_man_in_ff_w_lg_w_q_range146w148w(0) <= wire_man_in_ff_w_q_range146w(0) OR wire_w_man_not_zero_w_range144w(0);
	wire_man_in_ff_w_lg_w_q_range149w151w(0) <= wire_man_in_ff_w_q_range149w(0) OR wire_w_man_not_zero_w_range147w(0);
	wire_man_in_ff_w_lg_w_q_range152w154w(0) <= wire_man_in_ff_w_q_range152w(0) OR wire_w_man_not_zero_w_range150w(0);
	wire_man_in_ff_w_lg_w_q_range155w157w(0) <= wire_man_in_ff_w_q_range155w(0) OR wire_w_man_not_zero_w_range153w(0);
	wire_man_in_ff_w_lg_w_q_range158w160w(0) <= wire_man_in_ff_w_q_range158w(0) OR wire_w_man_not_zero_w_range156w(0);
	wire_man_in_ff_w_lg_w_q_range161w163w(0) <= wire_man_in_ff_w_q_range161w(0) OR wire_w_man_not_zero_w_range159w(0);
	wire_man_in_ff_w_lg_w_q_range164w166w(0) <= wire_man_in_ff_w_q_range164w(0) OR wire_w_man_not_zero_w_range162w(0);
	wire_man_in_ff_w_lg_w_q_range167w169w(0) <= wire_man_in_ff_w_q_range167w(0) OR wire_w_man_not_zero_w_range165w(0);
	wire_man_in_ff_w_lg_w_q_range170w172w(0) <= wire_man_in_ff_w_q_range170w(0) OR wire_w_man_not_zero_w_range168w(0);
	wire_man_in_ff_w_lg_w_q_range89w91w(0) <= wire_man_in_ff_w_q_range89w(0) OR wire_w_man_not_zero_w_range87w(0);
	wire_man_in_ff_w_lg_w_q_range173w175w(0) <= wire_man_in_ff_w_q_range173w(0) OR wire_w_man_not_zero_w_range171w(0);
	wire_man_in_ff_w_lg_w_q_range176w178w(0) <= wire_man_in_ff_w_q_range176w(0) OR wire_w_man_not_zero_w_range174w(0);
	wire_man_in_ff_w_lg_w_q_range179w181w(0) <= wire_man_in_ff_w_q_range179w(0) OR wire_w_man_not_zero_w_range177w(0);
	wire_man_in_ff_w_lg_w_q_range182w184w(0) <= wire_man_in_ff_w_q_range182w(0) OR wire_w_man_not_zero_w_range180w(0);
	wire_man_in_ff_w_lg_w_q_range185w187w(0) <= wire_man_in_ff_w_q_range185w(0) OR wire_w_man_not_zero_w_range183w(0);
	wire_man_in_ff_w_lg_w_q_range188w190w(0) <= wire_man_in_ff_w_q_range188w(0) OR wire_w_man_not_zero_w_range186w(0);
	wire_man_in_ff_w_lg_w_q_range191w193w(0) <= wire_man_in_ff_w_q_range191w(0) OR wire_w_man_not_zero_w_range189w(0);
	wire_man_in_ff_w_lg_w_q_range194w196w(0) <= wire_man_in_ff_w_q_range194w(0) OR wire_w_man_not_zero_w_range192w(0);
	wire_man_in_ff_w_lg_w_q_range197w199w(0) <= wire_man_in_ff_w_q_range197w(0) OR wire_w_man_not_zero_w_range195w(0);
	wire_man_in_ff_w_lg_w_q_range200w202w(0) <= wire_man_in_ff_w_q_range200w(0) OR wire_w_man_not_zero_w_range198w(0);
	wire_man_in_ff_w_lg_w_q_range92w94w(0) <= wire_man_in_ff_w_q_range92w(0) OR wire_w_man_not_zero_w_range90w(0);
	wire_man_in_ff_w_lg_w_q_range203w205w(0) <= wire_man_in_ff_w_q_range203w(0) OR wire_w_man_not_zero_w_range201w(0);
	wire_man_in_ff_w_lg_w_q_range206w208w(0) <= wire_man_in_ff_w_q_range206w(0) OR wire_w_man_not_zero_w_range204w(0);
	wire_man_in_ff_w_lg_w_q_range209w211w(0) <= wire_man_in_ff_w_q_range209w(0) OR wire_w_man_not_zero_w_range207w(0);
	wire_man_in_ff_w_lg_w_q_range212w214w(0) <= wire_man_in_ff_w_q_range212w(0) OR wire_w_man_not_zero_w_range210w(0);
	wire_man_in_ff_w_lg_w_q_range215w217w(0) <= wire_man_in_ff_w_q_range215w(0) OR wire_w_man_not_zero_w_range213w(0);
	wire_man_in_ff_w_lg_w_q_range218w220w(0) <= wire_man_in_ff_w_q_range218w(0) OR wire_w_man_not_zero_w_range216w(0);
	wire_man_in_ff_w_lg_w_q_range221w223w(0) <= wire_man_in_ff_w_q_range221w(0) OR wire_w_man_not_zero_w_range219w(0);
	wire_man_in_ff_w_lg_w_q_range224w226w(0) <= wire_man_in_ff_w_q_range224w(0) OR wire_w_man_not_zero_w_range222w(0);
	wire_man_in_ff_w_lg_w_q_range227w229w(0) <= wire_man_in_ff_w_q_range227w(0) OR wire_w_man_not_zero_w_range225w(0);
	wire_man_in_ff_w_lg_w_q_range230w232w(0) <= wire_man_in_ff_w_q_range230w(0) OR wire_w_man_not_zero_w_range228w(0);
	wire_man_in_ff_w_lg_w_q_range95w97w(0) <= wire_man_in_ff_w_q_range95w(0) OR wire_w_man_not_zero_w_range93w(0);
	wire_man_in_ff_w_lg_w_q_range233w235w(0) <= wire_man_in_ff_w_q_range233w(0) OR wire_w_man_not_zero_w_range231w(0);
	wire_man_in_ff_w_lg_w_q_range236w238w(0) <= wire_man_in_ff_w_q_range236w(0) OR wire_w_man_not_zero_w_range234w(0);
	wire_man_in_ff_w_lg_w_q_range98w100w(0) <= wire_man_in_ff_w_q_range98w(0) OR wire_w_man_not_zero_w_range96w(0);
	wire_man_in_ff_w_lg_w_q_range101w103w(0) <= wire_man_in_ff_w_q_range101w(0) OR wire_w_man_not_zero_w_range99w(0);
	wire_man_in_ff_w_lg_w_q_range104w106w(0) <= wire_man_in_ff_w_q_range104w(0) OR wire_w_man_not_zero_w_range102w(0);
	wire_man_in_ff_w_lg_w_q_range107w109w(0) <= wire_man_in_ff_w_q_range107w(0) OR wire_w_man_not_zero_w_range105w(0);
	wire_man_in_ff_w_lg_w_q_range110w112w(0) <= wire_man_in_ff_w_q_range110w(0) OR wire_w_man_not_zero_w_range108w(0);
	wire_man_in_ff_w_q_range83w(0) <= man_in_ff(0);
	wire_man_in_ff_w_q_range113w(0) <= man_in_ff(10);
	wire_man_in_ff_w_q_range116w(0) <= man_in_ff(11);
	wire_man_in_ff_w_q_range119w(0) <= man_in_ff(12);
	wire_man_in_ff_w_q_range122w(0) <= man_in_ff(13);
	wire_man_in_ff_w_q_range125w(0) <= man_in_ff(14);
	wire_man_in_ff_w_q_range128w(0) <= man_in_ff(15);
	wire_man_in_ff_w_q_range131w(0) <= man_in_ff(16);
	wire_man_in_ff_w_q_range134w(0) <= man_in_ff(17);
	wire_man_in_ff_w_q_range137w(0) <= man_in_ff(18);
	wire_man_in_ff_w_q_range140w(0) <= man_in_ff(19);
	wire_man_in_ff_w_q_range86w(0) <= man_in_ff(1);
	wire_man_in_ff_w_q_range143w(0) <= man_in_ff(20);
	wire_man_in_ff_w_q_range146w(0) <= man_in_ff(21);
	wire_man_in_ff_w_q_range149w(0) <= man_in_ff(22);
	wire_man_in_ff_w_q_range152w(0) <= man_in_ff(23);
	wire_man_in_ff_w_q_range155w(0) <= man_in_ff(24);
	wire_man_in_ff_w_q_range158w(0) <= man_in_ff(25);
	wire_man_in_ff_w_q_range161w(0) <= man_in_ff(26);
	wire_man_in_ff_w_q_range164w(0) <= man_in_ff(27);
	wire_man_in_ff_w_q_range167w(0) <= man_in_ff(28);
	wire_man_in_ff_w_q_range170w(0) <= man_in_ff(29);
	wire_man_in_ff_w_q_range89w(0) <= man_in_ff(2);
	wire_man_in_ff_w_q_range173w(0) <= man_in_ff(30);
	wire_man_in_ff_w_q_range176w(0) <= man_in_ff(31);
	wire_man_in_ff_w_q_range179w(0) <= man_in_ff(32);
	wire_man_in_ff_w_q_range182w(0) <= man_in_ff(33);
	wire_man_in_ff_w_q_range185w(0) <= man_in_ff(34);
	wire_man_in_ff_w_q_range188w(0) <= man_in_ff(35);
	wire_man_in_ff_w_q_range191w(0) <= man_in_ff(36);
	wire_man_in_ff_w_q_range194w(0) <= man_in_ff(37);
	wire_man_in_ff_w_q_range197w(0) <= man_in_ff(38);
	wire_man_in_ff_w_q_range200w(0) <= man_in_ff(39);
	wire_man_in_ff_w_q_range92w(0) <= man_in_ff(3);
	wire_man_in_ff_w_q_range203w(0) <= man_in_ff(40);
	wire_man_in_ff_w_q_range206w(0) <= man_in_ff(41);
	wire_man_in_ff_w_q_range209w(0) <= man_in_ff(42);
	wire_man_in_ff_w_q_range212w(0) <= man_in_ff(43);
	wire_man_in_ff_w_q_range215w(0) <= man_in_ff(44);
	wire_man_in_ff_w_q_range218w(0) <= man_in_ff(45);
	wire_man_in_ff_w_q_range221w(0) <= man_in_ff(46);
	wire_man_in_ff_w_q_range224w(0) <= man_in_ff(47);
	wire_man_in_ff_w_q_range227w(0) <= man_in_ff(48);
	wire_man_in_ff_w_q_range230w(0) <= man_in_ff(49);
	wire_man_in_ff_w_q_range95w(0) <= man_in_ff(4);
	wire_man_in_ff_w_q_range269w <= man_in_ff(50 DOWNTO 0);
	wire_man_in_ff_w_q_range233w(0) <= man_in_ff(50);
	wire_man_in_ff_w_q_range271w <= man_in_ff(51 DOWNTO 1);
	wire_man_in_ff_w_q_range236w(0) <= man_in_ff(51);
	wire_man_in_ff_w_q_range98w(0) <= man_in_ff(5);
	wire_man_in_ff_w_q_range101w(0) <= man_in_ff(6);
	wire_man_in_ff_w_q_range104w(0) <= man_in_ff(7);
	wire_man_in_ff_w_q_range107w(0) <= man_in_ff(8);
	wire_man_in_ff_w_q_range110w(0) <= man_in_ff(9);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_not_zero_ff <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_not_zero_ff <= man_not_zero_w(51);
			END IF;
		END IF;
	END PROCESS;
	wire_man_not_zero_ff_w_lg_q239w(0) <= NOT man_not_zero_ff;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_result_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_result_ff <= wire_man_rounding_ff_w_lg_w_lg_q285w286w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_rounding_ff <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_rounding_ff <= wire_add_sub3_result;
			END IF;
		END IF;
	END PROCESS;
	loop214 : FOR i IN 0 TO 51 GENERATE 
		wire_man_rounding_ff_w_lg_q285w(i) <= man_rounding_ff(i) AND zero_exp_ff26;
	END GENERATE loop214;
	loop215 : FOR i IN 0 TO 51 GENERATE 
		wire_man_rounding_ff_w_lg_w_lg_q285w286w(i) <= wire_man_rounding_ff_w_lg_q285w(i) OR nan_man_ff26;
	END GENERATE loop215;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff0 <= nancondition_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff1 <= nan_man_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff2 <= nan_man_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff3 <= nan_man_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff4 <= nan_man_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff5 <= nan_man_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff6 <= nan_man_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff7 <= nan_man_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff8 <= nan_man_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff9 <= nan_man_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff10 <= nan_man_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff11 <= nan_man_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff12 <= nan_man_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff13 <= nan_man_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff14 <= nan_man_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff15 <= nan_man_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff16 <= nan_man_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff17 <= nan_man_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff18 <= nan_man_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff19 <= nan_man_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff20 <= nan_man_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff21 <= nan_man_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff22 <= nan_man_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff23 <= nan_man_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff24 <= nan_man_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff25 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff25 <= nan_man_ff24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN nan_man_ff26 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN nan_man_ff26 <= nan_man_ff25;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff0 <= data(63);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff1 <= sign_node_ff0;
			END IF;
		END IF;
	END PROCESS;
	wire_sign_node_ff_w_lg_q244w(0) <= NOT sign_node_ff1;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff2 <= sign_node_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff3 <= sign_node_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff4 <= sign_node_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff5 <= sign_node_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff6 <= sign_node_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff7 <= sign_node_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff8 <= sign_node_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff9 <= sign_node_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff10 <= sign_node_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff11 <= sign_node_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff12 <= sign_node_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff13 <= sign_node_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff14 <= sign_node_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff15 <= sign_node_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff16 <= sign_node_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff17 <= sign_node_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff18 <= sign_node_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff19 <= sign_node_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff20 <= sign_node_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff21 <= sign_node_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff22 <= sign_node_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff23 <= sign_node_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff24 <= sign_node_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff25 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff25 <= sign_node_ff24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff26 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff26 <= sign_node_ff25;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff27 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff27 <= sign_node_ff26;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff28 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff28 <= sign_node_ff27;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_node_ff29 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_node_ff29 <= sign_node_ff28;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff0 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff0 <= exp_not_zero_ff;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff1 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff1 <= zero_exp_ff0;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff2 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff2 <= zero_exp_ff1;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff3 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff3 <= zero_exp_ff2;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff4 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff4 <= zero_exp_ff3;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff5 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff5 <= zero_exp_ff4;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff6 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff6 <= zero_exp_ff5;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff7 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff7 <= zero_exp_ff6;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff8 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff8 <= zero_exp_ff7;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff9 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff9 <= zero_exp_ff8;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff10 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff10 <= zero_exp_ff9;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff11 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff11 <= zero_exp_ff10;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff12 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff12 <= zero_exp_ff11;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff13 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff13 <= zero_exp_ff12;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff14 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff14 <= zero_exp_ff13;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff15 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff15 <= zero_exp_ff14;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff16 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff16 <= zero_exp_ff15;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff17 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff17 <= zero_exp_ff16;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff18 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff18 <= zero_exp_ff17;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff19 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff19 <= zero_exp_ff18;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff20 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff20 <= zero_exp_ff19;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff21 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff21 <= zero_exp_ff20;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff22 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff22 <= zero_exp_ff21;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff23 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff23 <= zero_exp_ff22;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff24 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff24 <= zero_exp_ff23;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff25 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff25 <= zero_exp_ff24;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN zero_exp_ff26 <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN zero_exp_ff26 <= zero_exp_ff25;
			END IF;
		END IF;
	END PROCESS;
	wire_add_sub1_dataa <= ( "0" & exp_in_ff);
	wire_add_sub1_datab <= ( "0" & bias);
	add_sub1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		dataa => wire_add_sub1_dataa,
		datab => wire_add_sub1_datab,
		result => wire_add_sub1_result
	  );
	wire_add_sub3_datab <= ( "000000000000000000000000000000000000000000000000000" & roundbit_w);
	add_sub3 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_PIPELINE => 0,
		LPM_WIDTH => 52
	  )
	  PORT MAP ( 
		dataa => man_root_result_w(52 DOWNTO 1),
		datab => wire_add_sub3_datab,
		result => wire_add_sub3_result
	  );

 END RTL; --fp_sqrt_dp_altfp_sqrt_lqd
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY fp_sqrt_dp IS
	PORT
	(
		aclr		: IN STD_LOGIC ;
		clk_en		: IN STD_LOGIC ;
		clock		: IN STD_LOGIC ;
		data		: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
END fp_sqrt_dp;


ARCHITECTURE RTL OF fp_sqrt_dp IS

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (63 DOWNTO 0);



	COMPONENT fp_sqrt_dp_altfp_sqrt_lqd
	PORT (
			clk_en	: IN STD_LOGIC ;
			clock	: IN STD_LOGIC ;
			aclr	: IN STD_LOGIC ;
			data	: IN STD_LOGIC_VECTOR (63 DOWNTO 0);
			result	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	result    <= sub_wire0(63 DOWNTO 0);

	fp_sqrt_dp_altfp_sqrt_lqd_component : fp_sqrt_dp_altfp_sqrt_lqd
	PORT MAP (
		clk_en => clk_en,
		clock => clock,
		aclr => aclr,
		data => data,
		result => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: FPM_FORMAT NUMERIC "1"
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Stratix II"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "30"
-- Retrieval info: CONSTANT: ROUNDING STRING "TO_NEAREST"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "11"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "52"
-- Retrieval info: USED_PORT: aclr 0 0 0 0 INPUT NODEFVAL "aclr"
-- Retrieval info: USED_PORT: clk_en 0 0 0 0 INPUT NODEFVAL "clk_en"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: data 0 0 64 0 INPUT NODEFVAL "data[63..0]"
-- Retrieval info: USED_PORT: result 0 0 64 0 OUTPUT NODEFVAL "result[63..0]"
-- Retrieval info: CONNECT: @data 0 0 64 0 data 0 0 64 0
-- Retrieval info: CONNECT: @clk_en 0 0 0 0 clk_en 0 0 0 0
-- Retrieval info: CONNECT: @aclr 0 0 0 0 aclr 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 64 0 @result 0 0 64 0
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_sqrt_dp.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_sqrt_dp.inc TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_sqrt_dp.cmp FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_sqrt_dp.bsf TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL fp_sqrt_dp_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
